* NGSPICE file created from Modulator.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

.subckt Modulator CLK_EXT CLK_PLL CLK_SR Data_SR NMOS1_PS1 NMOS1_PS2 NMOS2_PS1 NMOS2_PS2
+ NMOS_PS3 PMOS1_PS1 PMOS1_PS2 PMOS2_PS1 PMOS2_PS2 PMOS_PS3 RST SIGNAL_OUTPUT VGND
+ VPWR d1[0] d1[1] d1[2] d1[3] d1[4] d1[5] d2[0] d2[1] d2[2] d2[3] d2[4] d2[5]
XFILLER_0_27_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1270_ _0629_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_14_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0985_ _0443_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0770_ Signal_Generator_1_180phase_inst.count\[3\] Signal_Generator_1_180phase_inst.count\[2\]
+ _0284_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__and3_1
X_1253_ _0454_ _0455_ Dead_Time_Generator_inst_4.count_dt\[0\] VGND VGND VPWR VPWR
+ _0617_ sky130_fd_sc_hd__a21oi_1
X_1322_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0019_ _0105_ VGND VGND VPWR
+ VPWR Signal_Generator_1_270phase_inst.count\[5\] sky130_fd_sc_hd__dfstp_1
X_1184_ _0563_ _0564_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0968_ Shift_Register_Inst.data_out\[9\] Shift_Register_Inst.data_out\[10\] VGND
+ VGND VPWR VPWR _0430_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0899_ _0367_ _0378_ _0381_ Signal_Generator_2_180phase_inst.direction VGND VGND
+ VPWR VPWR _0038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0822_ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[1\]
+ Signal_Generator_2_0phase_inst.count\[3\] Signal_Generator_2_0phase_inst.count\[2\]
+ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__or4_2
XFILLER_0_28_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0753_ _0262_ _0269_ _0271_ Signal_Generator_1_90phase_inst.direction VGND VGND VPWR
+ VPWR _0023_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0684_ _0221_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__clkbuf_1
X_1305_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk net49 _0088_ VGND VGND VPWR
+ VPWR Signal_Generator_1_90phase_inst.count\[2\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_36_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1236_ _0603_ _0604_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1098_ _0499_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__inv_2
X_1167_ _0548_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__buf_2
XFILLER_0_40_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1021_ Shift_Register_Inst.data_out\[8\] Shift_Register_Inst.data_out\[7\] VGND VGND
+ VPWR VPWR _0460_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0805_ _0304_ _0309_ _0310_ Signal_Generator_1_270phase_inst.direction VGND VGND
+ VPWR VPWR _0015_ sky130_fd_sc_hd__a22o_1
X_0736_ Signal_Generator_1_0phase_inst.count\[4\] Signal_Generator_1_0phase_inst.direction
+ _0239_ Signal_Generator_1_0phase_inst.count\[5\] VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__o31a_1
XFILLER_0_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0667_ Shift_Register_Inst.shift_state\[1\] _0190_ _0196_ VGND VGND VPWR VPWR _0209_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_46_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1219_ Dead_Time_Generator_inst_2.count_dt\[3\] _0585_ Dead_Time_Generator_inst_2.count_dt\[4\]
+ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold52 Signal_Generator_2_90phase_inst.direction VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 Signal_Generator_2_180phase_inst.direction VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 Dead_Time_Generator_inst_1.count_dt\[4\] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1004_ _0441_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0719_ _0245_ _0242_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput20 net20 VGND VGND VPWR VPWR PMOS1_PS1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0984_ _0443_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1321_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0018_ _0104_ VGND VGND VPWR
+ VPWR Signal_Generator_1_270phase_inst.count\[4\] sky130_fd_sc_hd__dfrtp_4
X_1252_ Dead_Time_Generator_inst_4.count_dt\[0\] _0454_ _0455_ VGND VGND VPWR VPWR
+ _0616_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1183_ Dead_Time_Generator_inst_1.count_dt\[1\] net32 VGND VGND VPWR VPWR _0564_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_50 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0967_ net22 net20 net15 net17 _0428_ Shift_Register_Inst.data_out\[9\] VGND VGND
+ VPWR VPWR _0429_ sky130_fd_sc_hd__mux4_1
X_0898_ _0379_ _0380_ _0370_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0752_ net35 _0270_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0821_ Signal_Generator_1_270phase_inst.count\[4\] Signal_Generator_1_270phase_inst.direction
+ _0306_ _0322_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0683_ _0182_ Shift_Register_Inst.data_out\[9\] _0220_ VGND VGND VPWR VPWR _0221_
+ sky130_fd_sc_hd__mux2_1
X_1304_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0022_ _0087_ VGND VGND VPWR
+ VPWR Signal_Generator_1_90phase_inst.count\[1\] sky130_fd_sc_hd__dfstp_1
X_1235_ Dead_Time_Generator_inst_3.count_dt\[0\] _0603_ _0604_ VGND VGND VPWR VPWR
+ _0605_ sky130_fd_sc_hd__and3_1
X_1166_ _0514_ net45 _0542_ _0547_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__or4b_2
X_1097_ _0499_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__inv_2
X_1020_ Shift_Register_Inst.data_out\[7\] Shift_Register_Inst.data_out\[8\] VGND VGND
+ VPWR VPWR _0459_ sky130_fd_sc_hd__nor2b_2
XPHY_EDGE_ROW_28_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0735_ Signal_Generator_1_0phase_inst.direction _0256_ _0257_ _0241_ _0258_ VGND
+ VGND VPWR VPWR _0004_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_12_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0804_ _0307_ _0309_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__or2b_1
X_0666_ Shift_Register_Inst.data_out\[5\] VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__clkbuf_2
X_1218_ _0590_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
X_1149_ _0511_ _0512_ _0514_ _0530_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__o22a_1
Xhold53 Signal_Generator_1_0phase_inst.direction VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 _0546_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 Signal_Generator_2_270phase_inst.count\[0\] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 Dead_Time_Generator_inst_1.dt\[3\] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ _0444_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__inv_2
X_0718_ Signal_Generator_1_0phase_inst.count\[1\] Signal_Generator_1_0phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0649_ Shift_Register_Inst.shift_state\[0\] _0196_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__and2_1
Xoutput21 net21 VGND VGND VPWR VPWR PMOS1_PS2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_15_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0983_ _0443_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1320_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0017_ _0103_ VGND VGND VPWR
+ VPWR Signal_Generator_1_270phase_inst.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_1182_ Dead_Time_Generator_inst_1.count_dt\[1\] net32 VGND VGND VPWR VPWR _0563_
+ sky130_fd_sc_hd__nand2_1
X_1251_ _0615_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0897_ net65 Signal_Generator_2_180phase_inst.count\[1\] Signal_Generator_2_180phase_inst.count\[2\]
+ Signal_Generator_2_180phase_inst.count\[3\] VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__a31o_1
X_0966_ Shift_Register_Inst.data_out\[10\] VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0751_ Signal_Generator_1_90phase_inst.count\[2\] _0263_ VGND VGND VPWR VPWR _0270_
+ sky130_fd_sc_hd__xor2_1
X_0820_ Signal_Generator_1_270phase_inst.count\[4\] Signal_Generator_1_270phase_inst.direction
+ _0302_ Signal_Generator_1_270phase_inst.count\[5\] VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__o31a_1
XFILLER_0_3_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1303_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0021_ _0086_ VGND VGND VPWR
+ VPWR Signal_Generator_1_90phase_inst.count\[0\] sky130_fd_sc_hd__dfstp_1
X_0682_ _0188_ Shift_Register_Inst.shift_state\[2\] _0209_ VGND VGND VPWR VPWR _0220_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1096_ _0499_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__inv_2
X_1234_ net30 Dead_Time_Generator_inst_3.count_dt\[4\] VGND VGND VPWR VPWR _0604_
+ sky130_fd_sc_hd__or2b_1
X_1165_ _0529_ _0521_ _0528_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0949_ _0410_ _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0734_ Signal_Generator_1_0phase_inst.count\[4\] _0239_ VGND VGND VPWR VPWR _0258_
+ sky130_fd_sc_hd__xnor2_1
X_0665_ _0207_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0803_ _0308_ _0305_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__or2_1
X_1079_ _0498_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1148_ _0521_ _0528_ _0529_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__a21boi_1
X_1217_ _0545_ _0549_ _0589_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_45_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold10 _0265_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 Signal_Generator_1_180phase_inst.count\[0\] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 _0548_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 Dead_Time_Generator_inst_3.count_dt\[3\] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 Shift_Register_Inst.shift_state\[1\] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1002_ _0444_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0717_ net60 VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__inv_2
X_0648_ Shift_Register_Inst.shift_state\[1\] _0185_ net72 VGND VGND VPWR VPWR _0196_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput22 net22 VGND VGND VPWR VPWR PMOS2_PS1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0982_ _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1181_ _0545_ _0549_ net32 _0562_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__a211oi_1
X_1250_ _0544_ _0548_ _0614_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0896_ _0369_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__inv_2
X_0965_ Shift_Register_Inst.data_out\[12\] VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0750_ Signal_Generator_1_90phase_inst.count\[2\] net48 VGND VGND VPWR VPWR _0269_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0681_ _0219_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__clkbuf_1
X_1302_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk net36 _0085_ VGND VGND VPWR
+ VPWR Signal_Generator_1_90phase_inst.direction sky130_fd_sc_hd__dfstp_2
X_1233_ _0595_ net38 _0600_ _0601_ _0602_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__a221o_1
X_1095_ _0499_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__inv_2
X_1164_ _0522_ _0526_ _0527_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0948_ Dead_Time_Generator_inst_2.go net3 Shift_Register_Inst.data_out\[13\] VGND
+ VGND VPWR VPWR _0416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0879_ Signal_Generator_2_180phase_inst.direction VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0802_ Signal_Generator_1_270phase_inst.count\[1\] Signal_Generator_1_270phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__nor2_1
X_0733_ Signal_Generator_1_0phase_inst.count\[4\] _0243_ VGND VGND VPWR VPWR _0257_
+ sky130_fd_sc_hd__or2_1
X_0664_ _0182_ Dead_Time_Generator_inst_1.dt\[4\] _0206_ VGND VGND VPWR VPWR _0207_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1216_ _0569_ _0585_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__xnor2_1
X_1078_ _0441_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__buf_4
X_1147_ _0519_ _0520_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__nand2_1
Xhold11 _0027_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 Signal_Generator_1_90phase_inst.count\[1\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold44 _0173_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 Signal_Generator_1_270phase_inst.count\[0\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 Signal_Generator_1_270phase_inst.direction VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlygate4sd3_1
X_1001_ _0444_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_54 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0716_ _0241_ _0244_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0647_ _0192_ _0195_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput23 net23 VGND VGND VPWR VPWR PMOS2_PS2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0981_ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1180_ Dead_Time_Generator_inst_1.count_dt\[0\] _0561_ VGND VGND VPWR VPWR _0562_
+ sky130_fd_sc_hd__nor2_1
X_0964_ _0426_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
XFILLER_0_40_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0895_ _0365_ _0377_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0680_ _0182_ _0217_ _0218_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__mux2_1
X_1301_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0005_ _0084_ VGND VGND VPWR
+ VPWR Signal_Generator_1_0phase_inst.count\[5\] sky130_fd_sc_hd__dfrtp_2
X_1232_ Dead_Time_Generator_inst_3.count_dt\[4\] net64 VGND VGND VPWR VPWR _0602_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1094_ _0499_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__inv_2
X_1163_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__buf_2
X_0947_ _0415_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
XFILLER_0_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0878_ Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_180phase_inst.count\[1\]
+ Signal_Generator_2_180phase_inst.count\[3\] Signal_Generator_2_180phase_inst.count\[2\]
+ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__or4_2
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0801_ net58 VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__inv_2
X_0732_ _0253_ Signal_Generator_1_0phase_inst.count\[5\] Signal_Generator_1_0phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__or3b_1
X_0663_ _0183_ _0184_ _0193_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1215_ _0588_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__clkbuf_1
X_1146_ _0522_ _0526_ _0527_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__a21o_1
X_1077_ _0497_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold45 Signal_Generator_1_180phase_inst.direction VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 _0266_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 RST VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 Dead_Time_Generator_inst_3.count_dt\[4\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1000_ _0444_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0715_ Signal_Generator_1_0phase_inst.count\[5\] Signal_Generator_1_0phase_inst.count\[4\]
+ _0243_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__and3_1
X_0646_ _0189_ _0191_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1129_ _0510_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput24 net24 VGND VGND VPWR VPWR PMOS_PS3 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0980_ net2 VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_0__f_Dead_Time_Generator_inst_1.clk net26 VGND VGND VPWR VPWR clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_19_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0894_ net65 Signal_Generator_2_180phase_inst.count\[1\] Signal_Generator_2_180phase_inst.count\[2\]
+ Signal_Generator_2_180phase_inst.count\[3\] VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__o31ai_1
X_0963_ _0419_ _0423_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1300_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0004_ _0083_ VGND VGND VPWR
+ VPWR Signal_Generator_1_0phase_inst.count\[4\] sky130_fd_sc_hd__dfrtp_4
X_1162_ _0531_ _0542_ _0543_ _0539_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_0_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1231_ _0596_ Dead_Time_Generator_inst_1.dt\[2\] Dead_Time_Generator_inst_1.dt\[3\]
+ _0595_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1093_ _0499_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__inv_2
X_0877_ Signal_Generator_2_90phase_inst.count\[4\] Signal_Generator_2_90phase_inst.direction
+ _0348_ _0364_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__a31o_1
X_0946_ _0414_ _0410_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0731_ _0241_ _0252_ _0255_ Signal_Generator_1_0phase_inst.direction VGND VGND VPWR
+ VPWR _0003_ sky130_fd_sc_hd__a22o_1
X_0800_ _0304_ _0307_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__nor2_1
X_0662_ _0205_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1214_ _0545_ _0549_ _0587_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1145_ Shift_Register_Inst.data_out\[13\] net3 VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__or2b_1
X_1076_ _0497_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0929_ Signal_Generator_2_270phase_inst.count\[4\] _0390_ VGND VGND VPWR VPWR _0404_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_30_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold24 _0023_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 Signal_Generator_1_0phase_inst.count\[0\] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 Signal_Generator_2_90phase_inst.direction VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 Dead_Time_Generator_inst_1.dt\[3\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_7_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0714_ Signal_Generator_1_0phase_inst.count\[3\] Signal_Generator_1_0phase_inst.count\[2\]
+ _0242_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0645_ _0188_ _0192_ _0194_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__o21ai_1
X_1059_ _0445_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__inv_2
X_1128_ _0501_ _0502_ _0507_ _0508_ _0509_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__a32o_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput25 net25 VGND VGND VPWR VPWR SIGNAL_OUTPUT sky130_fd_sc_hd__buf_8
XFILLER_0_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0893_ _0367_ _0374_ _0376_ net66 VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__a22o_1
X_0962_ _0425_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
XFILLER_0_4_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1161_ net42 VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1092_ _0499_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__inv_2
X_1230_ _0596_ Dead_Time_Generator_inst_1.dt\[2\] _0597_ _0598_ _0599_ VGND VGND VPWR
+ VPWR _0600_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0876_ Signal_Generator_2_90phase_inst.count\[4\] Signal_Generator_2_90phase_inst.direction
+ _0344_ Signal_Generator_2_90phase_inst.count\[5\] VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__o31a_1
XFILLER_0_2_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0945_ _0413_ net4 Shift_Register_Inst.data_out\[13\] VGND VGND VPWR VPWR _0414_
+ sky130_fd_sc_hd__mux2_1
X_1359_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0166_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_2.count_dt\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0730_ _0253_ _0254_ _0244_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0661_ _0182_ Dead_Time_Generator_inst_1.dt\[3\] _0204_ VGND VGND VPWR VPWR _0205_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1213_ _0585_ _0586_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__nor2_1
X_1075_ _0497_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__inv_2
X_1144_ Signal_Generator_1_180phase_inst.count\[0\] _0503_ _0523_ _0524_ _0525_ VGND
+ VGND VPWR VPWR _0526_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_23_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0928_ _0400_ Signal_Generator_2_270phase_inst.count\[5\] Signal_Generator_2_270phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__or3b_1
X_0859_ _0350_ _0347_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold36 Signal_Generator_2_90phase_inst.count\[0\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 _0577_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 Dead_Time_Generator_inst_1.count_dt\[3\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 Shift_Register_Inst.shift_state\[4\] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0713_ Signal_Generator_1_0phase_inst.count\[1\] Signal_Generator_1_0phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__and2_1
X_0644_ _0191_ _0193_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1127_ Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[2\]
+ Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[2\]
+ Shift_Register_Inst.data_out\[5\] _0212_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__mux4_1
X_1058_ _0496_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput15 net15 VGND VGND VPWR VPWR NMOS1_PS1 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_25 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0961_ _0416_ _0421_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0892_ _0370_ _0375_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_56 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1160_ _0539_ _0540_ _0541_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__or3_1
X_1091_ _0499_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__inv_2
X_0944_ Dead_Time_Generator_inst_3.go VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0875_ net77 _0361_ _0362_ _0346_ _0363_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1358_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0165_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_2.count_dt\[1\] sky130_fd_sc_hd__dfxtp_1
X_1289_ clknet_1_1__leaf_CLK_SR _0152_ _0073_ VGND VGND VPWR VPWR Shift_Register_Inst.shift_state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0660_ _0185_ _0191_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1212_ Dead_Time_Generator_inst_2.count_dt\[1\] _0579_ Dead_Time_Generator_inst_2.count_dt\[2\]
+ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__a21oi_1
X_1074_ _0497_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__inv_2
X_1143_ _0208_ _0212_ Signal_Generator_1_270phase_inst.count\[0\] VGND VGND VPWR VPWR
+ _0525_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0927_ _0388_ _0399_ _0402_ Signal_Generator_2_270phase_inst.direction VGND VGND
+ VPWR VPWR _0045_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0789_ Signal_Generator_1_180phase_inst.count\[4\] _0285_ VGND VGND VPWR VPWR _0299_
+ sky130_fd_sc_hd__or2_1
X_0858_ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold37 Dead_Time_Generator_inst_3.count_dt\[0\] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 _0582_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 _0198_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 _0161_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0712_ Signal_Generator_1_0phase_inst.count\[5\] Signal_Generator_1_0phase_inst.count\[4\]
+ _0239_ _0240_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__o31a_2
X_0643_ _0188_ Shift_Register_Inst.shift_state\[2\] VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__nand2_1
X_1126_ Shift_Register_Inst.data_out\[13\] net5 VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__or2b_1
X_1057_ _0456_ _0492_ _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput16 net16 VGND VGND VPWR VPWR NMOS1_PS2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ _0500_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0960_ _0424_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_1
X_0891_ Signal_Generator_2_180phase_inst.count\[2\] _0368_ VGND VGND VPWR VPWR _0375_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1374_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0181_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_3.go sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1090_ _0499_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__inv_2
X_0874_ Signal_Generator_2_90phase_inst.count\[4\] _0344_ VGND VGND VPWR VPWR _0363_
+ sky130_fd_sc_hd__xnor2_1
X_0943_ _0412_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
XFILLER_0_27_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1357_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0164_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_2.count_dt\[0\] sky130_fd_sc_hd__dfxtp_1
X_1288_ clknet_1_1__leaf_CLK_SR _0151_ _0072_ VGND VGND VPWR VPWR Dead_Time_Generator_inst_1.dt\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1142_ Shift_Register_Inst.data_out\[6\] VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__inv_2
X_1211_ Dead_Time_Generator_inst_2.count_dt\[2\] Dead_Time_Generator_inst_2.count_dt\[1\]
+ _0579_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__and3_1
X_1073_ _0497_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__inv_2
X_0926_ _0400_ _0401_ _0391_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__a21o_1
X_0857_ net61 VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold38 Signal_Generator_1_90phase_inst.count\[0\] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlygate4sd3_1
X_0788_ _0295_ Signal_Generator_1_180phase_inst.count\[5\] Signal_Generator_1_180phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__or3b_1
Xhold27 Dead_Time_Generator_inst_1.count_dt\[2\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 Shift_Register_Inst.data_out\[16\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 Signal_Generator_1_180phase_inst.direction VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0711_ Signal_Generator_1_0phase_inst.direction VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_1__f_Dead_Time_Generator_inst_1.clk net26 VGND VGND VPWR VPWR clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk
+ sky130_fd_sc_hd__clkbuf_16
X_0642_ _0189_ _0191_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__nor2_1
X_1125_ Signal_Generator_1_180phase_inst.count\[3\] _0503_ _0504_ _0505_ _0506_ VGND
+ VGND VPWR VPWR _0507_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1056_ _0468_ _0480_ _0494_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__or3_1
Xoutput17 net17 VGND VGND VPWR VPWR NMOS2_PS1 sky130_fd_sc_hd__clkbuf_4
X_0909_ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1108_ _0500_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__inv_2
X_1039_ net12 _0470_ _0471_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_14 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0890_ Signal_Generator_2_180phase_inst.count\[2\] _0371_ VGND VGND VPWR VPWR _0374_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_2_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1373_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0180_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_4.count_dt\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0873_ Signal_Generator_2_90phase_inst.count\[4\] _0348_ VGND VGND VPWR VPWR _0362_
+ sky130_fd_sc_hd__or2_1
X_0942_ _0410_ _0411_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1356_ clknet_1_1__leaf_CLK_SR _0163_ _0134_ VGND VGND VPWR VPWR Dead_Time_Generator_inst_1.dt\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_1287_ clknet_1_1__leaf_CLK_SR _0150_ _0071_ VGND VGND VPWR VPWR Dead_Time_Generator_inst_1.dt\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1072_ _0497_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__inv_2
X_1141_ Signal_Generator_1_90phase_inst.count\[0\] _0208_ VGND VGND VPWR VPWR _0523_
+ sky130_fd_sc_hd__or2b_1
X_1210_ _0584_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0787_ _0283_ _0294_ _0297_ net70 VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__a22o_1
X_0856_ _0346_ _0349_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__nor2_1
X_0925_ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[1\]
+ Signal_Generator_2_270phase_inst.count\[2\] Signal_Generator_2_270phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold17 _0540_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 Dead_Time_Generator_inst_4.count_dt\[1\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 Dead_Time_Generator_inst_1.dt\[4\] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlygate4sd3_1
X_1339_ net29 _0036_ _0122_ VGND VGND VPWR VPWR Signal_Generator_2_180phase_inst.count\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_46_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0710_ Signal_Generator_1_0phase_inst.count\[3\] Signal_Generator_1_0phase_inst.count\[2\]
+ Signal_Generator_1_0phase_inst.count\[1\] Signal_Generator_1_0phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__or4_2
X_0641_ _0190_ _0183_ Shift_Register_Inst.shift_state\[1\] VGND VGND VPWR VPWR _0191_
+ sky130_fd_sc_hd__or3b_2
XFILLER_0_20_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1124_ net44 _0212_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_11_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1055_ _0486_ _0493_ _0489_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__or3b_1
X_0908_ Signal_Generator_2_270phase_inst.count\[5\] Signal_Generator_2_270phase_inst.count\[4\]
+ _0386_ _0387_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__o31a_1
Xoutput18 net18 VGND VGND VPWR VPWR NMOS2_PS2 sky130_fd_sc_hd__clkbuf_4
X_0839_ _0323_ _0335_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1107_ _0500_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__inv_2
X_1038_ _0472_ _0476_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1372_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0179_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_4.count_dt\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0941_ Dead_Time_Generator_inst_4.go net5 Shift_Register_Inst.data_out\[13\] VGND
+ VGND VPWR VPWR _0411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0872_ _0358_ Signal_Generator_2_90phase_inst.count\[5\] Signal_Generator_2_90phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__or3b_1
XFILLER_0_27_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1355_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0162_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_1.count_dt\[4\] sky130_fd_sc_hd__dfxtp_1
X_1286_ clknet_1_1__leaf_CLK_SR _0149_ _0070_ VGND VGND VPWR VPWR Dead_Time_Generator_inst_1.dt\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_41_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1071_ _0497_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__inv_2
X_1140_ _0000_ _0506_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0924_ _0390_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__inv_2
X_0786_ _0295_ _0296_ _0286_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__a21o_1
X_0855_ Signal_Generator_2_90phase_inst.count\[5\] Signal_Generator_2_90phase_inst.count\[4\]
+ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold18 _0159_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
X_1338_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0035_ _0121_ VGND VGND VPWR
+ VPWR Signal_Generator_2_180phase_inst.count\[0\] sky130_fd_sc_hd__dfstp_1
Xhold29 Signal_Generator_2_0phase_inst.count\[0\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
X_1269_ _0492_ _0495_ _0628_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0640_ Shift_Register_Inst.shift_state\[0\] VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1123_ Shift_Register_Inst.data_out\[5\] Shift_Register_Inst.data_out\[6\] Signal_Generator_1_270phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__and3_1
X_1054_ _0488_ _0487_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0907_ Signal_Generator_2_270phase_inst.direction VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0769_ Signal_Generator_1_180phase_inst.count\[1\] Signal_Generator_1_180phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__and2_1
Xoutput19 net19 VGND VGND VPWR VPWR NMOS_PS3 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0838_ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[1\]
+ Signal_Generator_2_0phase_inst.count\[2\] Signal_Generator_2_0phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__o31ai_1
XPHY_EDGE_ROW_44_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1106_ _0500_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__inv_2
X_1037_ _0474_ _0475_ net11 VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1371_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0178_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_4.count_dt\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0940_ Shift_Register_Inst.data_out\[15\] Shift_Register_Inst.data_out\[16\] Shift_Register_Inst.data_out\[17\]
+ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0871_ _0346_ _0357_ _0360_ net71 VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1285_ clknet_1_1__leaf_CLK_SR _0148_ _0069_ VGND VGND VPWR VPWR Dead_Time_Generator_inst_1.dt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1354_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk net51 VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_1.count_dt\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1070_ _0497_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__inv_2
X_0854_ Signal_Generator_2_90phase_inst.count\[3\] Signal_Generator_2_90phase_inst.count\[2\]
+ _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__and3_1
X_0923_ _0386_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__nand2_1
X_0785_ Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[1\]
+ Signal_Generator_1_180phase_inst.count\[0\] Signal_Generator_1_180phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold19 Shift_Register_Inst.data_out\[5\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1337_ net29 _0041_ _0120_ VGND VGND VPWR VPWR Signal_Generator_2_180phase_inst.direction
+ sky130_fd_sc_hd__dfstp_2
X_1268_ Dead_Time_Generator_inst_4.count_dt\[3\] _0622_ Dead_Time_Generator_inst_4.count_dt\[4\]
+ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__a21o_1
X_1199_ _0570_ Dead_Time_Generator_inst_1.dt\[2\] net38 _0569_ VGND VGND VPWR VPWR
+ _0575_ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1122_ Shift_Register_Inst.data_out\[6\] Signal_Generator_1_90phase_inst.count\[3\]
+ Shift_Register_Inst.data_out\[5\] VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__and3b_1
X_1053_ _0465_ _0466_ _0468_ _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_28_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0906_ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[1\]
+ Signal_Generator_2_270phase_inst.count\[3\] Signal_Generator_2_270phase_inst.count\[2\]
+ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__or4_2
X_0837_ _0325_ _0332_ _0334_ Signal_Generator_2_0phase_inst.direction VGND VGND VPWR
+ VPWR _0030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0768_ Signal_Generator_1_180phase_inst.count\[5\] Signal_Generator_1_180phase_inst.count\[4\]
+ _0281_ _0282_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__o31a_2
X_0699_ net1 Shift_Register_Inst.data_out\[14\] _0231_ VGND VGND VPWR VPWR _0232_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1105_ _0500_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1036_ Signal_Generator_2_0phase_inst.count\[2\] _0458_ VGND VGND VPWR VPWR _0475_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_16_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1019_ _0215_ _0217_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__nor2_2
XFILLER_0_8_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1370_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0177_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_4.count_dt\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_2__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VGND VPWR VPWR clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
X_0870_ _0358_ _0359_ _0349_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__a21o_1
X_1284_ clknet_1_1__leaf_CLK_SR _0147_ _0068_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_1353_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0160_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_1.count_dt\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0999_ _0444_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0922_ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[1\]
+ Signal_Generator_2_270phase_inst.count\[2\] Signal_Generator_2_270phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__o31ai_1
X_0853_ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0784_ _0285_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__inv_2
X_1336_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0054_ _0119_ VGND VGND VPWR
+ VPWR Signal_Generator_2_90phase_inst.count\[5\] sky130_fd_sc_hd__dfrtp_1
X_1267_ _0627_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__clkbuf_1
X_1198_ _0570_ Dead_Time_Generator_inst_1.dt\[2\] _0571_ _0572_ _0573_ VGND VGND VPWR
+ VPWR _0574_ sky130_fd_sc_hd__a221o_1
Xinput1 Data_SR VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
XFILLER_0_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1121_ Shift_Register_Inst.data_out\[5\] Shift_Register_Inst.data_out\[6\] VGND VGND
+ VPWR VPWR _0503_ sky130_fd_sc_hd__and2b_1
X_1052_ _0477_ _0478_ _0480_ _0490_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0767_ Signal_Generator_1_180phase_inst.direction VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__inv_2
X_0905_ Signal_Generator_2_180phase_inst.count\[4\] Signal_Generator_2_180phase_inst.direction
+ _0369_ _0385_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__a31o_1
X_0836_ _0328_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0698_ _0228_ _0201_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__or2_1
X_1319_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0016_ _0102_ VGND VGND VPWR
+ VPWR Signal_Generator_1_270phase_inst.count\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1035_ Signal_Generator_2_180phase_inst.count\[2\] _0459_ _0460_ Signal_Generator_2_90phase_inst.count\[2\]
+ _0473_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__a221oi_2
X_1104_ _0500_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0819_ Signal_Generator_1_270phase_inst.direction _0319_ _0320_ _0304_ _0321_ VGND
+ VGND VPWR VPWR _0018_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1018_ _0215_ _0217_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1283_ clknet_1_1__leaf_CLK_SR _0146_ _0067_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_1352_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk net43 VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_1.count_dt\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0998_ _0444_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0921_ _0388_ _0395_ _0397_ Signal_Generator_2_270phase_inst.direction VGND VGND
+ VPWR VPWR _0044_ sky130_fd_sc_hd__a22o_1
X_0783_ _0281_ _0293_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__nand2_1
X_0852_ Signal_Generator_2_90phase_inst.count\[5\] Signal_Generator_2_90phase_inst.count\[4\]
+ _0344_ _0345_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__o31a_2
XFILLER_0_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1335_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0053_ _0118_ VGND VGND VPWR
+ VPWR Signal_Generator_2_90phase_inst.count\[4\] sky130_fd_sc_hd__dfstp_2
Xinput2 net37 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1266_ _0593_ _0594_ _0626_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__and3_1
X_1197_ Dead_Time_Generator_inst_2.count_dt\[1\] Dead_Time_Generator_inst_1.dt\[1\]
+ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1120_ _0208_ _0212_ Signal_Generator_1_0phase_inst.count\[3\] VGND VGND VPWR VPWR
+ _0502_ sky130_fd_sc_hd__or3_1
X_1051_ _0486_ _0489_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0904_ Signal_Generator_2_180phase_inst.count\[4\] Signal_Generator_2_180phase_inst.direction
+ _0365_ Signal_Generator_2_180phase_inst.count\[5\] VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__o31a_1
XFILLER_0_28_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0766_ Signal_Generator_1_180phase_inst.count\[3\] Signal_Generator_1_180phase_inst.count\[2\]
+ Signal_Generator_1_180phase_inst.count\[1\] Signal_Generator_1_180phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__or4_2
X_0835_ Signal_Generator_2_0phase_inst.count\[2\] _0326_ VGND VGND VPWR VPWR _0333_
+ sky130_fd_sc_hd__xor2_1
X_0697_ _0230_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1318_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0015_ _0101_ VGND VGND VPWR
+ VPWR Signal_Generator_1_270phase_inst.count\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1249_ _0577_ _0578_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1103_ _0500_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__inv_2
X_1034_ _0215_ _0217_ Signal_Generator_2_270phase_inst.count\[2\] VGND VGND VPWR VPWR
+ _0473_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0749_ _0262_ _0267_ _0268_ Signal_Generator_1_90phase_inst.direction VGND VGND VPWR
+ VPWR _0022_ sky130_fd_sc_hd__a22o_1
X_0818_ Signal_Generator_1_270phase_inst.count\[4\] _0302_ VGND VGND VPWR VPWR _0321_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1017_ _0454_ _0455_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1351_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk net33 VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_1.count_dt\[0\] sky130_fd_sc_hd__dfxtp_1
X_1282_ clknet_1_1__leaf_CLK_SR _0145_ _0066_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0997_ _0444_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0920_ _0391_ _0396_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__or2_1
X_0782_ Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[1\]
+ Signal_Generator_1_180phase_inst.count\[0\] Signal_Generator_1_180phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__o31ai_1
X_0851_ Signal_Generator_2_90phase_inst.direction VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__inv_2
X_1334_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0052_ _0117_ VGND VGND VPWR
+ VPWR Signal_Generator_2_90phase_inst.count\[3\] sky130_fd_sc_hd__dfstp_1
X_1265_ _0446_ _0622_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 d1[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
X_1196_ Dead_Time_Generator_inst_2.count_dt\[0\] Dead_Time_Generator_inst_1.dt\[0\]
+ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1050_ net10 _0485_ _0487_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_43_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0903_ Signal_Generator_2_180phase_inst.direction _0382_ _0383_ _0367_ _0384_ VGND
+ VGND VPWR VPWR _0039_ sky130_fd_sc_hd__a32o_1
X_0834_ Signal_Generator_2_0phase_inst.count\[2\] _0329_ VGND VGND VPWR VPWR _0332_
+ sky130_fd_sc_hd__xor2_1
X_0765_ Signal_Generator_1_90phase_inst.count\[4\] Signal_Generator_1_90phase_inst.direction
+ _0264_ _0280_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0696_ net1 Shift_Register_Inst.data_out\[13\] _0229_ VGND VGND VPWR VPWR _0230_
+ sky130_fd_sc_hd__mux2_1
X_1248_ _0593_ _0594_ _0612_ net59 VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__o2bb2a_1
X_1317_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0014_ _0100_ VGND VGND VPWR
+ VPWR Signal_Generator_1_270phase_inst.count\[0\] sky130_fd_sc_hd__dfrtp_2
X_1179_ _0558_ net31 VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1102_ _0500_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1033_ _0470_ _0471_ net12 VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_16_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0817_ Signal_Generator_1_270phase_inst.count\[4\] _0306_ VGND VGND VPWR VPWR _0320_
+ sky130_fd_sc_hd__or2_1
X_0748_ _0265_ _0267_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__or2b_1
X_0679_ _0183_ _0188_ Shift_Register_Inst.shift_state\[2\] _0184_ VGND VGND VPWR VPWR
+ _0218_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_39_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1016_ net30 Dead_Time_Generator_inst_4.count_dt\[4\] VGND VGND VPWR VPWR _0455_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1350_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0047_ _0133_ VGND VGND VPWR
+ VPWR Signal_Generator_2_270phase_inst.count\[5\] sky130_fd_sc_hd__dfstp_1
X_1281_ clknet_1_0__leaf_CLK_SR _0144_ _0065_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0996_ _0444_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0850_ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[1\]
+ Signal_Generator_2_90phase_inst.count\[3\] Signal_Generator_2_90phase_inst.count\[2\]
+ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__or4_2
X_0781_ _0283_ _0290_ _0292_ net70 VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1333_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0051_ _0116_ VGND VGND VPWR
+ VPWR Signal_Generator_2_90phase_inst.count\[2\] sky130_fd_sc_hd__dfstp_2
X_1264_ _0625_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__clkbuf_1
Xinput4 d1[1] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1195_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_2.count_dt\[1\]
+ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__or2b_1
X_0979_ _0427_ _0434_ _0440_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__a21bo_4
XFILLER_0_43_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0902_ Signal_Generator_2_180phase_inst.count\[4\] _0365_ VGND VGND VPWR VPWR _0384_
+ sky130_fd_sc_hd__xnor2_1
X_0833_ _0325_ _0330_ _0331_ Signal_Generator_2_0phase_inst.direction VGND VGND VPWR
+ VPWR _0029_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0764_ Signal_Generator_1_90phase_inst.count\[4\] Signal_Generator_1_90phase_inst.direction
+ _0260_ Signal_Generator_1_90phase_inst.count\[5\] VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__o31a_1
X_0695_ _0228_ _0209_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__or2_1
X_1247_ _0593_ _0594_ _0612_ _0613_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__a211oi_1
X_1316_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0020_ _0099_ VGND VGND VPWR
+ VPWR Signal_Generator_1_270phase_inst.direction sky130_fd_sc_hd__dfrtp_4
X_1178_ Dead_Time_Generator_inst_1.count_dt\[0\] _0558_ net31 VGND VGND VPWR VPWR
+ _0560_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1101_ _0500_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__inv_2
X_1032_ Signal_Generator_2_0phase_inst.count\[3\] _0458_ VGND VGND VPWR VPWR _0471_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0747_ _0266_ _0263_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__or2_1
X_0816_ _0316_ Signal_Generator_1_270phase_inst.count\[5\] Signal_Generator_1_270phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__or3b_1
XFILLER_0_42_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0678_ Shift_Register_Inst.data_out\[8\] VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_39_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_3__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VGND VPWR VPWR clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1015_ _0446_ net38 _0451_ _0452_ _0453_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1280_ clknet_1_0__leaf_CLK_SR _0143_ _0064_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_0995_ _0444_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0780_ _0286_ _0291_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1332_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0050_ _0115_ VGND VGND VPWR
+ VPWR Signal_Generator_2_90phase_inst.count\[1\] sky130_fd_sc_hd__dfstp_1
X_1263_ _0593_ _0594_ _0624_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__and3_1
Xinput5 d1[2] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
X_1194_ Dead_Time_Generator_inst_2.count_dt\[2\] VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0978_ Shift_Register_Inst.data_out\[11\] _0427_ _0436_ _0439_ Shift_Register_Inst.data_out\[9\]
+ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__o32a_2
XFILLER_0_37_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0763_ Signal_Generator_1_90phase_inst.direction _0277_ _0278_ _0262_ _0279_ VGND
+ VGND VPWR VPWR _0025_ sky130_fd_sc_hd__a32o_1
X_0901_ Signal_Generator_2_180phase_inst.count\[4\] _0369_ VGND VGND VPWR VPWR _0383_
+ sky130_fd_sc_hd__or2_1
X_0832_ _0328_ _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__or2b_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1315_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0012_ _0098_ VGND VGND VPWR
+ VPWR Signal_Generator_1_180phase_inst.count\[5\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0694_ Shift_Register_Inst.shift_state\[3\] Shift_Register_Inst.shift_state\[2\]
+ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__nand2_1
X_1246_ _0596_ _0608_ _0595_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__o21a_1
X_1177_ net30 Dead_Time_Generator_inst_1.count_dt\[4\] VGND VGND VPWR VPWR _0559_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1031_ Signal_Generator_2_180phase_inst.count\[3\] _0459_ _0460_ Signal_Generator_2_90phase_inst.count\[3\]
+ _0469_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__a221oi_2
X_1100_ _0441_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0746_ net47 Signal_Generator_1_90phase_inst.count\[0\] VGND VGND VPWR VPWR _0266_
+ sky130_fd_sc_hd__nor2_1
X_0815_ _0304_ _0315_ _0318_ net80 VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0677_ _0216_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__clkbuf_1
X_1229_ Dead_Time_Generator_inst_3.count_dt\[1\] Dead_Time_Generator_inst_1.dt\[1\]
+ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_7_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ Dead_Time_Generator_inst_4.count_dt\[4\] Dead_Time_Generator_inst_1.dt\[4\]
+ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0729_ Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[1\]
+ Signal_Generator_1_0phase_inst.count\[0\] Signal_Generator_1_0phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0994_ _0444_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_39_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1331_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0049_ _0114_ VGND VGND VPWR
+ VPWR Signal_Generator_2_90phase_inst.count\[0\] sky130_fd_sc_hd__dfstp_1
X_1262_ _0622_ _0623_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__nor2_1
Xinput6 d1[3] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
X_1193_ Dead_Time_Generator_inst_2.count_dt\[3\] VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0977_ _0438_ Shift_Register_Inst.data_out\[10\] VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__nand2_2
XFILLER_0_37_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_194 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0379_ Signal_Generator_2_180phase_inst.count\[5\] Signal_Generator_2_180phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__or3b_1
X_0762_ Signal_Generator_1_90phase_inst.count\[4\] _0260_ VGND VGND VPWR VPWR _0279_
+ sky130_fd_sc_hd__xnor2_1
X_0831_ _0329_ _0326_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__or2_1
X_0693_ _0227_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1314_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0011_ _0097_ VGND VGND VPWR
+ VPWR Signal_Generator_1_180phase_inst.count\[4\] sky130_fd_sc_hd__dfstp_2
Xclkbuf_0_Dead_Time_Generator_inst_1.clk Dead_Time_Generator_inst_1.clk VGND VGND
+ VPWR VPWR clknet_0_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
X_1245_ Dead_Time_Generator_inst_3.count_dt\[3\] Dead_Time_Generator_inst_3.count_dt\[2\]
+ Dead_Time_Generator_inst_3.count_dt\[1\] _0605_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_19_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1176_ _0550_ net67 _0555_ _0556_ _0557_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1030_ _0215_ _0217_ Signal_Generator_2_270phase_inst.count\[3\] VGND VGND VPWR VPWR
+ _0469_ sky130_fd_sc_hd__and3_1
X_0814_ _0316_ _0317_ _0307_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0745_ net63 VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_10_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0676_ _0182_ _0215_ _0194_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1228_ Dead_Time_Generator_inst_3.count_dt\[0\] Dead_Time_Generator_inst_1.dt\[0\]
+ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__and2b_1
X_1159_ _0532_ _0533_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_7_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1013_ _0447_ Dead_Time_Generator_inst_1.dt\[2\] Dead_Time_Generator_inst_1.dt\[3\]
+ _0446_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0728_ _0243_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0659_ _0203_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_41_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0993_ _0441_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1330_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0055_ _0113_ VGND VGND VPWR
+ VPWR Signal_Generator_2_90phase_inst.direction sky130_fd_sc_hd__dfstp_1
X_1261_ net53 _0616_ Dead_Time_Generator_inst_4.count_dt\[2\] VGND VGND VPWR VPWR
+ _0623_ sky130_fd_sc_hd__a21oi_1
Xinput7 d1[4] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
X_1192_ _0442_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0976_ Shift_Register_Inst.data_out\[11\] _0427_ net23 _0437_ VGND VGND VPWR VPWR
+ _0438_ sky130_fd_sc_hd__a31o_4
XFILLER_0_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0830_ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__nor2_1
X_0761_ Signal_Generator_1_90phase_inst.count\[4\] _0264_ VGND VGND VPWR VPWR _0278_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_11_138 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0692_ net1 Shift_Register_Inst.data_out\[12\] _0226_ VGND VGND VPWR VPWR _0227_
+ sky130_fd_sc_hd__mux2_1
X_1313_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0010_ _0096_ VGND VGND VPWR
+ VPWR Signal_Generator_1_180phase_inst.count\[3\] sky130_fd_sc_hd__dfstp_1
X_1244_ _0593_ _0594_ _0611_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_19_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1175_ Dead_Time_Generator_inst_1.count_dt\[4\] net30 VGND VGND VPWR VPWR _0557_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0959_ _0414_ _0423_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0813_ Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[1\]
+ Signal_Generator_1_270phase_inst.count\[0\] Signal_Generator_1_270phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__a31o_1
Xinput10 d2[1] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
X_0744_ _0262_ net35 VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__nor2_1
X_0675_ Shift_Register_Inst.data_out\[7\] VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__clkbuf_2
X_1227_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_3.count_dt\[1\]
+ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__or2b_1
X_1158_ _0534_ _0538_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__nor2_1
X_1089_ _0441_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__buf_4
XFILLER_0_30_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1012_ _0447_ Dead_Time_Generator_inst_1.dt\[2\] _0448_ _0449_ _0450_ VGND VGND VPWR
+ VPWR _0451_ sky130_fd_sc_hd__a221o_1
X_0727_ _0239_ _0251_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__nand2_1
X_0658_ _0182_ Dead_Time_Generator_inst_1.dt\[2\] _0202_ VGND VGND VPWR VPWR _0203_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0992_ _0443_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput8 d1[5] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
X_1260_ Dead_Time_Generator_inst_4.count_dt\[2\] Dead_Time_Generator_inst_4.count_dt\[1\]
+ _0616_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__and3_1
X_1191_ _0545_ _0549_ _0567_ net55 VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__o2bb2a_1
X_0975_ Shift_Register_Inst.data_out\[11\] Shift_Register_Inst.data_out\[12\] clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__and3b_2
XFILLER_0_45_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_4__f_Dead_Time_Generator_inst_1.clk net28 VGND VGND VPWR VPWR clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0760_ _0274_ Signal_Generator_1_90phase_inst.count\[5\] Signal_Generator_1_90phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__or3b_1
XFILLER_0_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_47 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0691_ _0183_ _0188_ _0189_ _0184_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__or4_1
X_1312_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0009_ _0095_ VGND VGND VPWR
+ VPWR Signal_Generator_1_180phase_inst.count\[2\] sky130_fd_sc_hd__dfstp_2
X_1243_ _0596_ _0608_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__xnor2_1
X_1174_ _0551_ Dead_Time_Generator_inst_1.dt\[2\] Dead_Time_Generator_inst_1.dt\[3\]
+ _0550_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_19_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0889_ _0367_ _0372_ _0373_ Signal_Generator_2_180phase_inst.direction VGND VGND
+ VPWR VPWR _0036_ sky130_fd_sc_hd__a22o_1
X_0958_ Shift_Register_Inst.data_out\[16\] Shift_Register_Inst.data_out\[17\] Shift_Register_Inst.data_out\[15\]
+ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0743_ net34 Signal_Generator_1_90phase_inst.count\[4\] _0264_ VGND VGND VPWR VPWR
+ _0265_ sky130_fd_sc_hd__and3_1
X_0812_ _0306_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__inv_2
Xinput11 d2[2] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
XFILLER_0_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0674_ _0214_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__clkbuf_1
X_1157_ _0532_ _0533_ _0534_ _0538_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__a22o_1
X_1226_ net75 VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__inv_2
X_1088_ _0498_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1011_ Dead_Time_Generator_inst_4.count_dt\[1\] Dead_Time_Generator_inst_1.dt\[1\]
+ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__and2b_1
X_0726_ Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[1\]
+ Signal_Generator_1_0phase_inst.count\[0\] Signal_Generator_1_0phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_4_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0657_ _0185_ _0201_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__or2_1
X_1209_ _0545_ _0549_ _0583_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0709_ _0238_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_46_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0991_ _0443_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_46 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 d2[0] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_1190_ _0545_ _0549_ _0567_ _0568_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0974_ net24 _0430_ _0435_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0690_ _0225_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1311_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0008_ _0094_ VGND VGND VPWR
+ VPWR Signal_Generator_1_180phase_inst.count\[1\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1242_ _0593_ _0594_ _0610_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1173_ _0551_ Dead_Time_Generator_inst_1.dt\[2\] _0552_ _0553_ _0554_ VGND VGND VPWR
+ VPWR _0555_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_19_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0888_ _0370_ _0372_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__or2b_1
X_0957_ _0422_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
XFILLER_0_18_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0742_ Signal_Generator_1_90phase_inst.count\[3\] Signal_Generator_1_90phase_inst.count\[2\]
+ _0263_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__and3_1
X_0811_ _0302_ _0314_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__nand2_1
X_0673_ _0182_ _0212_ _0213_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__mux2_1
Xinput12 d2[3] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1156_ Signal_Generator_1_0phase_inst.count\[5\] _0506_ _0535_ _0537_ VGND VGND VPWR
+ VPWR _0538_ sky130_fd_sc_hd__a211o_1
X_1087_ _0498_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__inv_2
X_1225_ net68 VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1010_ Dead_Time_Generator_inst_4.count_dt\[0\] Dead_Time_Generator_inst_1.dt\[0\]
+ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_44_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0725_ _0241_ _0248_ _0250_ net78 VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__a22o_1
X_0656_ _0183_ Shift_Register_Inst.shift_state\[0\] Shift_Register_Inst.shift_state\[1\]
+ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_4_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1208_ Dead_Time_Generator_inst_2.count_dt\[1\] _0579_ VGND VGND VPWR VPWR _0583_
+ sky130_fd_sc_hd__xor2_1
X_1139_ _0519_ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0639_ Shift_Register_Inst.shift_state\[2\] VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__inv_2
X_0708_ net1 Shift_Register_Inst.data_out\[17\] _0237_ VGND VGND VPWR VPWR _0238_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0990_ _0443_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_17_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0973_ Shift_Register_Inst.data_out\[9\] _0428_ net19 VGND VGND VPWR VPWR _0435_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_2_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1310_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0007_ _0093_ VGND VGND VPWR
+ VPWR Signal_Generator_1_180phase_inst.count\[0\] sky130_fd_sc_hd__dfstp_2
X_1241_ _0608_ _0609_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1172_ Dead_Time_Generator_inst_1.count_dt\[1\] Dead_Time_Generator_inst_1.dt\[1\]
+ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0956_ _0411_ _0421_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0887_ _0371_ _0368_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0810_ Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[1\]
+ Signal_Generator_1_270phase_inst.count\[0\] Signal_Generator_1_270phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__o31ai_1
Xinput13 d2[4] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
X_0741_ net47 Signal_Generator_1_90phase_inst.count\[0\] VGND VGND VPWR VPWR _0263_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0672_ _0193_ _0201_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__or2_1
X_1224_ _0495_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__buf_2
X_1155_ Signal_Generator_1_180phase_inst.count\[5\] _0503_ _0536_ VGND VGND VPWR VPWR
+ _0537_ sky130_fd_sc_hd__a21o_1
X_1086_ _0498_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0939_ Shift_Register_Inst.data_out\[16\] _0409_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_38_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0724_ _0244_ _0249_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0655_ _0200_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_4_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1207_ net40 VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkbuf_1
X_1069_ _0497_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__inv_2
X_1138_ Shift_Register_Inst.data_out\[13\] net4 VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_31_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0707_ Shift_Register_Inst.shift_state\[1\] _0190_ _0185_ _0183_ VGND VGND VPWR VPWR
+ _0237_ sky130_fd_sc_hd__or4b_1
X_0638_ Shift_Register_Inst.shift_state\[3\] VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0972_ _0429_ _0433_ Shift_Register_Inst.data_out\[11\] VGND VGND VPWR VPWR _0434_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1240_ Dead_Time_Generator_inst_3.count_dt\[1\] _0605_ VGND VGND VPWR VPWR _0609_
+ sky130_fd_sc_hd__or2_1
X_1171_ Dead_Time_Generator_inst_1.count_dt\[0\] Dead_Time_Generator_inst_1.dt\[0\]
+ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0886_ net65 Signal_Generator_2_180phase_inst.count\[1\] VGND VGND VPWR VPWR _0371_
+ sky130_fd_sc_hd__nor2_1
X_0955_ Shift_Register_Inst.data_out\[16\] Shift_Register_Inst.data_out\[17\] Shift_Register_Inst.data_out\[15\]
+ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__and3b_1
XFILLER_0_27_231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1369_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0176_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_4.count_dt\[0\] sky130_fd_sc_hd__dfxtp_1
X_0740_ net34 Signal_Generator_1_90phase_inst.count\[4\] _0260_ _0261_ VGND VGND VPWR
+ VPWR _0262_ sky130_fd_sc_hd__o31a_1
Xinput14 d2[5] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
X_0671_ Shift_Register_Inst.data_out\[6\] VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1154_ Shift_Register_Inst.data_out\[5\] Shift_Register_Inst.data_out\[6\] Signal_Generator_1_270phase_inst.count\[5\]
+ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__and3_1
X_1223_ _0492_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__buf_2
X_1085_ _0498_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__inv_2
X_0869_ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[1\]
+ Signal_Generator_2_90phase_inst.count\[2\] Signal_Generator_2_90phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0938_ net7 VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0723_ Signal_Generator_1_0phase_inst.count\[2\] _0242_ VGND VGND VPWR VPWR _0249_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0654_ _0182_ Dead_Time_Generator_inst_1.dt\[1\] _0199_ VGND VGND VPWR VPWR _0200_
+ sky130_fd_sc_hd__mux2_1
X_1137_ _0506_ _0515_ _0516_ _0517_ _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__o41a_1
X_1206_ _0545_ _0549_ _0581_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__and3_1
X_1068_ _0497_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0706_ _0236_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_5__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VGND VPWR VPWR clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
X_0637_ net76 Shift_Register_Inst.shift_state\[2\] Shift_Register_Inst.shift_state\[1\]
+ Shift_Register_Inst.shift_state\[0\] _0183_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_0_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0971_ net21 _0430_ _0431_ net16 _0432_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_1.count_dt\[1\]
+ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__or2b_1
X_0885_ net65 VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__inv_2
X_0954_ _0420_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
XFILLER_0_27_243 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1299_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0003_ _0082_ VGND VGND VPWR
+ VPWR Signal_Generator_1_0phase_inst.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_1368_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0175_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_2.go sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0670_ _0211_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__clkbuf_1
X_1153_ _0208_ _0524_ Signal_Generator_1_90phase_inst.count\[5\] VGND VGND VPWR VPWR
+ _0535_ sky130_fd_sc_hd__and3_1
X_1084_ _0498_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__inv_2
X_1222_ _0545_ _0549_ _0561_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0868_ _0348_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__inv_2
X_0937_ _0408_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlymetal6s2s_1
X_0799_ Signal_Generator_1_270phase_inst.count\[5\] Signal_Generator_1_270phase_inst.count\[4\]
+ _0306_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0722_ Signal_Generator_1_0phase_inst.count\[2\] _0245_ VGND VGND VPWR VPWR _0248_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0653_ _0183_ Shift_Register_Inst.shift_state\[1\] _0190_ _0185_ VGND VGND VPWR VPWR
+ _0199_ sky130_fd_sc_hd__or4_1
X_1067_ _0441_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__buf_4
X_1136_ _0208_ _0212_ Signal_Generator_1_0phase_inst.count\[1\] VGND VGND VPWR VPWR
+ _0518_ sky130_fd_sc_hd__or3_1
X_1205_ _0579_ _0580_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0636_ _0187_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
X_0705_ net1 Shift_Register_Inst.data_out\[16\] _0235_ VGND VGND VPWR VPWR _0236_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1119_ Shift_Register_Inst.data_out\[13\] net6 VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0970_ Shift_Register_Inst.data_out\[9\] _0428_ net18 VGND VGND VPWR VPWR _0432_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0884_ _0367_ _0370_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0953_ _0419_ _0410_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__or2b_1
XFILLER_0_27_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1367_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0174_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_3.count_dt\[4\] sky130_fd_sc_hd__dfxtp_1
X_1298_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0002_ _0081_ VGND VGND VPWR
+ VPWR Signal_Generator_1_0phase_inst.count\[2\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_18_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1221_ _0592_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f_CLK_SR clknet_0_CLK_SR VGND VGND VPWR VPWR clknet_1_1__leaf_CLK_SR
+ sky130_fd_sc_hd__clkbuf_16
X_1083_ _0498_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__inv_2
X_1152_ net41 net8 VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__or2b_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0936_ Shift_Register_Inst.data_out\[16\] net8 VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__and2_1
X_0867_ _0344_ _0356_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0798_ Signal_Generator_1_270phase_inst.count\[3\] Signal_Generator_1_270phase_inst.count\[2\]
+ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0721_ _0241_ _0246_ _0247_ Signal_Generator_1_0phase_inst.direction VGND VGND VPWR
+ VPWR _0001_ sky130_fd_sc_hd__a22o_1
X_0652_ _0197_ net73 VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1204_ net39 _0578_ Dead_Time_Generator_inst_2.count_dt\[0\] VGND VGND VPWR VPWR
+ _0580_ sky130_fd_sc_hd__a21oi_1
X_1066_ _0445_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__inv_2
X_1135_ _0208_ _0212_ Signal_Generator_1_270phase_inst.count\[1\] VGND VGND VPWR VPWR
+ _0517_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_35_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0919_ Signal_Generator_2_270phase_inst.count\[2\] _0389_ VGND VGND VPWR VPWR _0396_
+ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_9_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 Dead_Time_Generator_inst_1.dt\[4\] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0635_ _0182_ Dead_Time_Generator_inst_1.dt\[0\] _0186_ VGND VGND VPWR VPWR _0187_
+ sky130_fd_sc_hd__mux2_1
X_0704_ Shift_Register_Inst.shift_state\[1\] Shift_Register_Inst.shift_state\[0\]
+ _0185_ _0183_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_0_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1118_ _0442_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__inv_2
X_1049_ net9 VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_23_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0952_ _0418_ net6 Shift_Register_Inst.data_out\[13\] VGND VGND VPWR VPWR _0419_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0883_ Signal_Generator_2_180phase_inst.count\[5\] Signal_Generator_2_180phase_inst.count\[4\]
+ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1366_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk net69 VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_3.count_dt\[3\] sky130_fd_sc_hd__dfxtp_1
X_1297_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0001_ _0080_ VGND VGND VPWR
+ VPWR Signal_Generator_1_0phase_inst.count\[1\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_18_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1151_ Signal_Generator_1_0phase_inst.count\[4\] Signal_Generator_1_90phase_inst.count\[4\]
+ Signal_Generator_1_180phase_inst.count\[4\] Signal_Generator_1_270phase_inst.count\[4\]
+ _0208_ _0212_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__mux4_1
X_1220_ _0544_ net46 _0591_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__and3_1
X_1082_ _0498_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__inv_2
X_0866_ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[1\]
+ Signal_Generator_2_90phase_inst.count\[2\] Signal_Generator_2_90phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_15_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0935_ _0407_ VGND VGND VPWR VPWR Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__buf_6
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0797_ Signal_Generator_1_270phase_inst.count\[1\] Signal_Generator_1_270phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__and2_1
X_1349_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0046_ _0132_ VGND VGND VPWR
+ VPWR Signal_Generator_2_270phase_inst.count\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0720_ _0244_ _0246_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_12_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0651_ Shift_Register_Inst.shift_state\[0\] _0196_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__nor2_1
X_1134_ _0212_ Signal_Generator_1_90phase_inst.count\[1\] _0208_ VGND VGND VPWR VPWR
+ _0516_ sky130_fd_sc_hd__and3b_1
XFILLER_0_18_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1203_ Dead_Time_Generator_inst_2.count_dt\[0\] _0577_ _0578_ VGND VGND VPWR VPWR
+ _0579_ sky130_fd_sc_hd__and3_1
X_1065_ _0445_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_35_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0918_ Signal_Generator_2_270phase_inst.count\[2\] _0392_ VGND VGND VPWR VPWR _0395_
+ sky130_fd_sc_hd__xor2_1
X_0849_ Signal_Generator_2_0phase_inst.count\[4\] Signal_Generator_2_0phase_inst.direction
+ _0327_ _0343_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold6 _0559_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_40_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0703_ _0234_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__clkbuf_1
X_0634_ _0183_ _0184_ _0185_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__or3_1
XFILLER_0_29_84 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1117_ _0442_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1048_ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[0\]
+ Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[0\]
+ _0215_ _0217_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_23_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0882_ Signal_Generator_2_180phase_inst.count\[3\] Signal_Generator_2_180phase_inst.count\[2\]
+ _0368_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0951_ Dead_Time_Generator_inst_1.go VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1296_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0000_ _0079_ VGND VGND VPWR
+ VPWR Signal_Generator_1_0phase_inst.count\[0\] sky130_fd_sc_hd__dfrtp_1
X_1365_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0172_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_3.count_dt\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1150_ net41 _0409_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__or2_1
X_1081_ _0498_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__inv_2
Xclkbuf_3_6__f_Dead_Time_Generator_inst_1.clk net27 VGND VGND VPWR VPWR clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
+ sky130_fd_sc_hd__clkbuf_16
X_0865_ _0346_ _0353_ _0355_ net71 VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__a22o_1
X_0934_ CLK_PLL CLK_EXT Shift_Register_Inst.data_out\[14\] VGND VGND VPWR VPWR _0407_
+ sky130_fd_sc_hd__mux2_4
X_0796_ Signal_Generator_1_270phase_inst.count\[5\] Signal_Generator_1_270phase_inst.count\[4\]
+ _0302_ _0303_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__o31a_1
X_1348_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0045_ _0131_ VGND VGND VPWR
+ VPWR Signal_Generator_2_270phase_inst.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_1279_ clknet_1_0__leaf_CLK_SR _0142_ _0063_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0650_ net79 _0197_ _0191_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__o21a_1
X_1064_ _0445_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__inv_2
X_1133_ _0208_ _0212_ Signal_Generator_1_180phase_inst.count\[1\] VGND VGND VPWR VPWR
+ _0515_ sky130_fd_sc_hd__and3b_1
XFILLER_0_18_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1202_ net30 Dead_Time_Generator_inst_2.count_dt\[4\] VGND VGND VPWR VPWR _0578_
+ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_35_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0779_ Signal_Generator_1_180phase_inst.count\[2\] _0284_ VGND VGND VPWR VPWR _0291_
+ sky130_fd_sc_hd__xor2_1
X_0917_ _0388_ _0393_ _0394_ Signal_Generator_2_270phase_inst.direction VGND VGND
+ VPWR VPWR _0043_ sky130_fd_sc_hd__a22o_1
X_0848_ Signal_Generator_2_0phase_inst.count\[4\] Signal_Generator_2_0phase_inst.direction
+ _0323_ Signal_Generator_2_0phase_inst.count\[5\] VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_3_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_CLK_SR CLK_SR VGND VGND VPWR VPWR clknet_0_CLK_SR sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold7 _0560_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
XFILLER_0_44_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0702_ net1 Shift_Register_Inst.data_out\[15\] _0233_ VGND VGND VPWR VPWR _0234_
+ sky130_fd_sc_hd__mux2_1
X_0633_ Shift_Register_Inst.shift_state\[3\] Shift_Register_Inst.shift_state\[2\]
+ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__or2_2
XFILLER_0_45_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1116_ _0442_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__inv_2
X_1047_ net10 _0485_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_87 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0881_ Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_180phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__and2_1
X_0950_ _0417_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
XFILLER_0_27_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1295_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0006_ _0078_ VGND VGND VPWR
+ VPWR Signal_Generator_1_0phase_inst.direction sky130_fd_sc_hd__dfstp_2
X_1364_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0171_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_3.count_dt\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1080_ _0498_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0795_ Signal_Generator_1_270phase_inst.direction VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__inv_2
X_0864_ _0349_ _0354_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__or2_1
X_0933_ Signal_Generator_2_270phase_inst.count\[4\] Signal_Generator_2_270phase_inst.direction
+ _0390_ _0406_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__a31o_1
X_1347_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0044_ _0130_ VGND VGND VPWR
+ VPWR Signal_Generator_2_270phase_inst.count\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1278_ clknet_1_0__leaf_CLK_SR _0141_ _0062_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_12_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1201_ _0569_ net38 _0574_ _0575_ _0576_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__a221o_1
X_1063_ _0445_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1132_ _0510_ _0512_ _0513_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_43_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0916_ _0391_ _0393_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__or2b_1
X_0778_ Signal_Generator_1_180phase_inst.count\[2\] _0287_ VGND VGND VPWR VPWR _0290_
+ sky130_fd_sc_hd__xor2_1
X_0847_ Signal_Generator_2_0phase_inst.direction _0340_ _0341_ _0325_ _0342_ VGND
+ VGND VPWR VPWR _0032_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_3_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 _0158_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0701_ _0228_ _0191_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__or2_1
X_0632_ Shift_Register_Inst.shift_state\[1\] Shift_Register_Inst.shift_state\[0\]
+ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1115_ _0442_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__inv_2
X_1046_ _0458_ _0481_ _0482_ _0483_ _0484_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__o41ai_1
XFILLER_0_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1029_ _0466_ _0467_ _0465_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__or3b_1
XFILLER_0_16_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0880_ Signal_Generator_2_180phase_inst.count\[5\] Signal_Generator_2_180phase_inst.count\[4\]
+ _0365_ _0366_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__o31a_2
XFILLER_0_12_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1363_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0170_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_3.count_dt\[0\] sky130_fd_sc_hd__dfxtp_1
X_1294_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0157_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_4.go sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0932_ Signal_Generator_2_270phase_inst.count\[4\] Signal_Generator_2_270phase_inst.direction
+ _0386_ Signal_Generator_2_270phase_inst.count\[5\] VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__o31a_1
XFILLER_0_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0794_ Signal_Generator_1_270phase_inst.count\[3\] Signal_Generator_1_270phase_inst.count\[2\]
+ Signal_Generator_1_270phase_inst.count\[1\] Signal_Generator_1_270phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__or4_2
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0863_ Signal_Generator_2_90phase_inst.count\[2\] _0347_ VGND VGND VPWR VPWR _0354_
+ sky130_fd_sc_hd__xor2_1
X_1346_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0043_ _0129_ VGND VGND VPWR
+ VPWR Signal_Generator_2_270phase_inst.count\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1277_ clknet_1_1__leaf_CLK_SR _0140_ _0061_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1200_ Dead_Time_Generator_inst_2.count_dt\[4\] net30 VGND VGND VPWR VPWR _0576_
+ sky130_fd_sc_hd__and2b_1
X_1062_ _0445_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__inv_2
X_1131_ _0508_ _0509_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_43_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0915_ _0392_ _0389_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__or2_1
X_0777_ _0283_ _0288_ _0289_ net70 VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0846_ Signal_Generator_2_0phase_inst.count\[4\] _0323_ VGND VGND VPWR VPWR _0342_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1329_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0033_ _0112_ VGND VGND VPWR
+ VPWR Signal_Generator_2_0phase_inst.count\[5\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_26_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 Signal_Generator_1_90phase_inst.count\[5\] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
X_0700_ _0232_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_29_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0631_ Shift_Register_Inst.shift_state\[4\] VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__clkbuf_2
X_1114_ _0442_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1045_ _0215_ _0217_ Signal_Generator_2_0phase_inst.count\[1\] VGND VGND VPWR VPWR
+ _0484_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0829_ net54 VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1028_ net13 _0464_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1362_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0169_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_1.go sky130_fd_sc_hd__dfxtp_1
X_1293_ clknet_1_1__leaf_CLK_SR _0156_ _0077_ VGND VGND VPWR VPWR Shift_Register_Inst.shift_state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0931_ Signal_Generator_2_270phase_inst.direction _0403_ _0404_ _0388_ _0405_ VGND
+ VGND VPWR VPWR _0046_ sky130_fd_sc_hd__a32o_1
X_0862_ Signal_Generator_2_90phase_inst.count\[2\] _0350_ VGND VGND VPWR VPWR _0353_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_15_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0793_ Signal_Generator_1_180phase_inst.count\[4\] Signal_Generator_1_180phase_inst.direction
+ _0285_ _0301_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__a31o_1
Xrebuffer1 clknet_0_Dead_Time_Generator_inst_1.clk VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_8
X_1345_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0042_ _0128_ VGND VGND VPWR
+ VPWR Signal_Generator_2_270phase_inst.count\[0\] sky130_fd_sc_hd__dfrtp_2
X_1276_ clknet_1_0__leaf_CLK_SR _0139_ _0060_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_38_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1130_ _0502_ _0507_ _0501_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1061_ _0445_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0914_ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__nor2_1
X_0845_ Signal_Generator_2_0phase_inst.count\[4\] _0327_ VGND VGND VPWR VPWR _0341_
+ sky130_fd_sc_hd__or2_1
X_0776_ _0286_ _0288_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__or2b_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1259_ _0621_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__clkbuf_1
X_1328_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0032_ _0111_ VGND VGND VPWR
+ VPWR Signal_Generator_2_0phase_inst.count\[4\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_26_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0630_ net1 VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__buf_2
XFILLER_0_29_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1044_ _0215_ _0217_ Signal_Generator_2_270phase_inst.count\[1\] VGND VGND VPWR VPWR
+ _0483_ sky130_fd_sc_hd__and3_1
X_1113_ _0442_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__inv_2
X_0759_ _0262_ _0273_ _0276_ Signal_Generator_1_90phase_inst.direction VGND VGND VPWR
+ VPWR _0024_ sky130_fd_sc_hd__a22o_1
X_0828_ _0325_ _0328_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_46_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1027_ net14 _0462_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_7__f_Dead_Time_Generator_inst_1.clk net27 VGND VGND VPWR VPWR clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1292_ clknet_1_1__leaf_CLK_SR _0155_ _0076_ VGND VGND VPWR VPWR Shift_Register_Inst.shift_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1361_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0168_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_2.count_dt\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0792_ Signal_Generator_1_180phase_inst.count\[4\] Signal_Generator_1_180phase_inst.direction
+ _0281_ Signal_Generator_1_180phase_inst.count\[5\] VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__o31a_1
X_0861_ _0346_ _0351_ _0352_ net71 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__a22o_1
X_0930_ Signal_Generator_2_270phase_inst.count\[4\] _0386_ VGND VGND VPWR VPWR _0405_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_15_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer2 clknet_0_Dead_Time_Generator_inst_1.clk VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1344_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0048_ _0127_ VGND VGND VPWR
+ VPWR Signal_Generator_2_270phase_inst.direction sky130_fd_sc_hd__dfrtp_4
X_1275_ clknet_1_0__leaf_CLK_SR _0138_ _0059_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1060_ _0445_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0775_ _0287_ _0284_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__or2_1
X_0913_ net56 VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__inv_2
X_0844_ _0337_ Signal_Generator_2_0phase_inst.count\[5\] Signal_Generator_2_0phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__or3b_1
X_1258_ _0593_ _0594_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__and3_1
X_1327_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0031_ _0110_ VGND VGND VPWR
+ VPWR Signal_Generator_2_0phase_inst.count\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1189_ _0551_ _0563_ _0550_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1112_ _0442_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__inv_2
X_1043_ _0215_ _0217_ Signal_Generator_2_180phase_inst.count\[1\] VGND VGND VPWR VPWR
+ _0482_ sky130_fd_sc_hd__and3b_1
XFILLER_0_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0758_ _0274_ _0275_ _0265_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0827_ Signal_Generator_2_0phase_inst.count\[5\] Signal_Generator_2_0phase_inst.count\[4\]
+ _0327_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__and3_1
X_0689_ net1 Shift_Register_Inst.data_out\[11\] _0224_ VGND VGND VPWR VPWR _0225_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1026_ net14 _0462_ _0464_ net13 VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__o22a_1
XFILLER_0_39_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1009_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_4.count_dt\[1\]
+ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__or2b_1
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1360_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0167_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_2.count_dt\[3\] sky130_fd_sc_hd__dfxtp_1
X_1291_ clknet_1_0__leaf_CLK_SR _0154_ _0075_ VGND VGND VPWR VPWR Shift_Register_Inst.shift_state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0791_ net74 _0298_ _0299_ _0283_ _0300_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__a32o_1
X_0860_ _0349_ _0351_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__or2b_1
Xrebuffer3 clknet_0_Dead_Time_Generator_inst_1.clk VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd1_1
X_1343_ net29 _0040_ _0126_ VGND VGND VPWR VPWR Signal_Generator_2_180phase_inst.count\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1274_ clknet_1_0__leaf_CLK_SR _0137_ _0058_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0989_ _0443_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0912_ _0388_ _0391_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__nor2_1
X_0774_ Signal_Generator_1_180phase_inst.count\[1\] Signal_Generator_1_180phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0843_ _0325_ _0336_ _0339_ Signal_Generator_2_0phase_inst.direction VGND VGND VPWR
+ VPWR _0031_ sky130_fd_sc_hd__a22o_1
X_1326_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0030_ _0109_ VGND VGND VPWR
+ VPWR Signal_Generator_2_0phase_inst.count\[2\] sky130_fd_sc_hd__dfrtp_4
X_1257_ Dead_Time_Generator_inst_4.count_dt\[1\] _0616_ VGND VGND VPWR VPWR _0620_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_26_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1188_ Dead_Time_Generator_inst_1.count_dt\[3\] Dead_Time_Generator_inst_1.count_dt\[2\]
+ Dead_Time_Generator_inst_1.count_dt\[1\] net32 VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__and4_1
XFILLER_0_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1111_ _0442_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__inv_2
X_1042_ _0217_ Signal_Generator_2_90phase_inst.count\[1\] _0215_ VGND VGND VPWR VPWR
+ _0481_ sky130_fd_sc_hd__and3b_1
XFILLER_0_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0757_ Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[1\]
+ Signal_Generator_1_90phase_inst.count\[0\] Signal_Generator_1_90phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__a31o_1
X_0826_ Signal_Generator_2_0phase_inst.count\[3\] Signal_Generator_2_0phase_inst.count\[2\]
+ _0326_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__and3_1
X_0688_ _0188_ Shift_Register_Inst.shift_state\[2\] _0191_ VGND VGND VPWR VPWR _0224_
+ sky130_fd_sc_hd__or3_1
X_1309_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0013_ _0092_ VGND VGND VPWR
+ VPWR Signal_Generator_1_180phase_inst.direction sky130_fd_sc_hd__dfstp_1
XFILLER_0_43_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1025_ Signal_Generator_2_270phase_inst.count\[4\] _0457_ _0458_ Signal_Generator_2_0phase_inst.count\[4\]
+ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__a221oi_2
X_0809_ _0304_ _0311_ _0313_ Signal_Generator_1_270phase_inst.direction VGND VGND
+ VPWR VPWR _0016_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1008_ Dead_Time_Generator_inst_4.count_dt\[2\] VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1290_ clknet_1_1__leaf_CLK_SR _0153_ _0074_ VGND VGND VPWR VPWR Shift_Register_Inst.shift_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0790_ Signal_Generator_1_180phase_inst.count\[4\] _0281_ VGND VGND VPWR VPWR _0300_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer4 clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk VGND VGND VPWR VPWR net29
+ sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1342_ net29 _0039_ _0125_ VGND VGND VPWR VPWR Signal_Generator_2_180phase_inst.count\[4\]
+ sky130_fd_sc_hd__dfstp_2
X_1273_ clknet_1_0__leaf_CLK_SR _0136_ _0057_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_0988_ _0443_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0911_ Signal_Generator_2_270phase_inst.count\[5\] Signal_Generator_2_270phase_inst.count\[4\]
+ _0390_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__and3_1
X_0842_ _0337_ _0338_ _0328_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__a21o_1
X_0773_ net57 VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1256_ _0619_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__clkbuf_1
X_1325_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0029_ _0108_ VGND VGND VPWR
+ VPWR Signal_Generator_2_0phase_inst.count\[1\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_34_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1187_ _0545_ _0549_ _0566_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1110_ _0500_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1041_ _0472_ _0476_ _0478_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__or4_1
X_0825_ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0756_ _0264_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__inv_2
X_0687_ _0223_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__clkbuf_1
X_1308_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0026_ _0091_ VGND VGND VPWR
+ VPWR Signal_Generator_1_90phase_inst.count\[5\] sky130_fd_sc_hd__dfrtp_1
X_1239_ Dead_Time_Generator_inst_3.count_dt\[1\] _0605_ VGND VGND VPWR VPWR _0608_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1024_ Signal_Generator_2_180phase_inst.count\[4\] _0459_ _0460_ Signal_Generator_2_90phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__a22o_1
X_0808_ _0307_ _0312_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__or2_1
X_0739_ Signal_Generator_1_90phase_inst.direction VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1007_ Dead_Time_Generator_inst_4.count_dt\[3\] VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_CLK_SR clknet_0_CLK_SR VGND VGND VPWR VPWR clknet_1_0__leaf_CLK_SR
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_44_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1341_ net29 _0038_ _0124_ VGND VGND VPWR VPWR Signal_Generator_2_180phase_inst.count\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1272_ clknet_1_0__leaf_CLK_SR _0135_ _0056_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0987_ _0443_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0772_ _0283_ _0286_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__nor2_1
X_0910_ Signal_Generator_2_270phase_inst.count\[3\] Signal_Generator_2_270phase_inst.count\[2\]
+ _0389_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_11_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0841_ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[1\]
+ Signal_Generator_2_0phase_inst.count\[2\] Signal_Generator_2_0phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1324_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0028_ _0107_ VGND VGND VPWR
+ VPWR Signal_Generator_2_0phase_inst.count\[0\] sky130_fd_sc_hd__dfrtp_2
X_1255_ _0593_ _0594_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__and3_1
X_1186_ _0551_ _0563_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_34_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1040_ net11 _0474_ _0475_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0755_ _0260_ _0272_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__nand2_1
X_0824_ Signal_Generator_2_0phase_inst.count\[5\] Signal_Generator_2_0phase_inst.count\[4\]
+ _0323_ _0324_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__o31a_2
XPHY_EDGE_ROW_24_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0686_ net1 Shift_Register_Inst.data_out\[10\] _0222_ VGND VGND VPWR VPWR _0223_
+ sky130_fd_sc_hd__mux2_1
X_1307_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0025_ _0090_ VGND VGND VPWR
+ VPWR Signal_Generator_1_90phase_inst.count\[4\] sky130_fd_sc_hd__dfstp_2
X_1238_ _0593_ _0594_ _0605_ _0607_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__a211oi_1
X_1169_ net52 VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1023_ Signal_Generator_2_270phase_inst.count\[5\] _0457_ _0458_ Signal_Generator_2_0phase_inst.count\[5\]
+ _0461_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__a221oi_2
X_0738_ Signal_Generator_1_90phase_inst.count\[3\] Signal_Generator_1_90phase_inst.count\[2\]
+ Signal_Generator_1_90phase_inst.count\[1\] Signal_Generator_1_90phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__or4_2
X_0807_ Signal_Generator_1_270phase_inst.count\[2\] _0305_ VGND VGND VPWR VPWR _0312_
+ sky130_fd_sc_hd__xor2_1
X_0669_ _0182_ _0208_ _0210_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 Dead_Time_Generator_inst_3.count_dt\[2\] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1006_ _0445_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1340_ net29 _0037_ _0123_ VGND VGND VPWR VPWR Signal_Generator_2_180phase_inst.count\[2\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_23_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1271_ _0593_ _0594_ _0606_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0986_ _0443_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0771_ Signal_Generator_1_180phase_inst.count\[5\] Signal_Generator_1_180phase_inst.count\[4\]
+ _0285_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__and3_1
X_0840_ _0327_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__inv_2
X_1323_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0034_ _0106_ VGND VGND VPWR
+ VPWR Signal_Generator_2_0phase_inst.direction sky130_fd_sc_hd__dfstp_2
X_1254_ _0616_ _0617_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__nor2_1
X_1185_ _0545_ _0549_ _0565_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0969_ Shift_Register_Inst.data_out\[9\] Shift_Register_Inst.data_out\[10\] VGND
+ VGND VPWR VPWR _0431_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0754_ Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[1\]
+ Signal_Generator_1_90phase_inst.count\[0\] Signal_Generator_1_90phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__o31ai_1
X_0823_ Signal_Generator_2_0phase_inst.direction VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__inv_2
X_0685_ _0188_ Shift_Register_Inst.shift_state\[2\] _0201_ VGND VGND VPWR VPWR _0222_
+ sky130_fd_sc_hd__or3_1
X_1306_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0024_ _0089_ VGND VGND VPWR
+ VPWR Signal_Generator_1_90phase_inst.count\[3\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_19_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1099_ _0499_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__inv_2
X_1237_ net62 _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__nor2_1
X_1168_ net50 VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1022_ Signal_Generator_2_180phase_inst.count\[5\] _0459_ _0460_ Signal_Generator_2_90phase_inst.count\[5\]
+ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0737_ Signal_Generator_1_0phase_inst.count\[4\] Signal_Generator_1_0phase_inst.direction
+ _0243_ _0259_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__a31o_1
X_0806_ Signal_Generator_1_270phase_inst.count\[2\] _0308_ VGND VGND VPWR VPWR _0311_
+ sky130_fd_sc_hd__xor2_1
X_0668_ _0193_ _0209_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold40 Signal_Generator_2_180phase_inst.count\[0\] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold51 Shift_Register_Inst.shift_state\[3\] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1005_ _0445_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

