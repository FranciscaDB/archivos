* NGSPICE file created from Modulator.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.226 ps=2.26 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.143 ps=1.62 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B X C VGND VPWR VNB VPB
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_4 VGND VPWR X B1 A2 A1 A3 VNB VPB
X0 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5 a_277_47# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_193_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_361_47# A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VGND A3 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X15 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X16 a_277_47# A1 a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_445_47# A2 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.5 pd=3 as=0.135 ps=1.27 w=1 l=0.15
X22 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X23 a_277_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.226 ps=2.26 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.143 ps=1.62 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR X A3 A2 A1 B1 B2 VNB VPB
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_2 VPWR VGND Q SET_B D CLK VNB VPB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X3 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X5 a_1228_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X6 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X8 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X10 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X11 VPWR a_1602_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1028_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VGND a_1602_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1028_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X20 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X21 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0441 ps=0.63 w=0.42 l=0.15
X23 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.223 pd=2.21 as=0.121 ps=1.16 w=0.84 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_1300_47# a_1178_261# a_1228_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X29 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X30 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X31 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.121 pd=1.16 as=0.109 ps=1.36 w=0.42 l=0.15
X32 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X33 VGND SET_B a_1300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0441 ps=0.63 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_1 VGND VPWR C B A Y VNB VPB
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_4 VGND VPWR A1 A2 B2 Y B1 VNB VPB
X0 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X17 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X30 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X31 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.226 ps=2.26 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.143 ps=1.62 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VNB VPB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 VPWR VGND A X B VNB VPB
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.226 ps=2.26 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.143 ps=1.62 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__a21o_1 VPWR VGND A2 A1 B1 X VNB VPB
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 VGND VPWR A B Y VNB VPB
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR X A1 S A0 VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 VPWR VGND Y A VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND B1 A1 A2 X B2 VNB VPB
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND B C A X VNB VPB
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 X A VGND VPWR VNB VPB
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR A X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_4 VGND VPWR X A B C VNB VPB
X0 VPWR A a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.198 pd=1.39 as=0.305 ps=2.61 w=1 l=0.15
X1 a_294_47# B a_185_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.128 ps=1.04 w=0.65 l=0.15
X2 a_185_47# A a_94_47# VNB sky130_fd_pr__nfet_01v8 ad=0.128 pd=1.04 as=0.198 ps=1.91 w=0.65 l=0.15
X3 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND C a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.08 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_94_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.198 ps=1.39 w=1 l=0.15
X6 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.177 ps=1.36 w=1 l=0.15
X7 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR C a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.36 as=0.14 ps=1.28 w=1 l=0.15
X9 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138 ps=1.08 w=0.65 l=0.15
X10 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_1 VPWR VGND Q SET_B D CLK VNB VPB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X6 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.123 ps=1.17 w=0.84 l=0.15
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 X A3 A2 A1 B1 VGND VPWR VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 VGND VPWR B C_N A X VNB VPB
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.1 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 Q CLK D VPWR VGND VNB VPB
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_1 VGND VPWR X A1 A2 B1 C1 VNB VPB
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 X A1 A2 A3 B1 VGND VPWR VNB VPB
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.213 ps=1.42 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_1 VGND VPWR A X B_N VNB VPB
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.157 ps=1.17 w=0.42 l=0.15
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 VGND VPWR A1 A2 B1 X VNB VPB
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 VGND VPWR X A2 B1 A1 C1 VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_2 VPWR VGND A2 A1 Y B1 C1 VNB VPB
X0 VGND A2 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR A1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_37_297# B1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_485_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_292_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VPWR A2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_485_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X11 a_37_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 Y A1 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X13 Y C1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14 a_292_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15 a_292_297# B1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND A2 A1 B1 Y VNB VPB
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X B A C VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR A X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 VGND VPWR CLK D RESET_B Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 VGND VPWR X A B VNB VPB
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 VGND VPWR B2 A2 A1 B1 X VNB VPB
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 VGND VPWR CLK D RESET_B Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_1 VPWR VGND X A1 A2 A3 B2 B1 VNB VPB
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.127 ps=1.04 w=0.65 l=0.15
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.133 ps=1.06 w=0.65 l=0.15
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.107 ps=0.98 w=0.65 l=0.15
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_2 VPWR VGND B D C A X VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.91 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 VGND VPWR A Y B VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 B1 Y A1 VNB VPB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND X A VNB VPB
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 Y B1 VPWR VGND VNB VPB
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.198 ps=1.26 w=0.65 l=0.15
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.393 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.393 ps=1.78 w=1 l=0.15
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 VGND VPWR B1 A1_N A2_N X B2 VNB VPB
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VGND VPWR A X VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR B Y A VNB VPB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_8 VGND VPWR A X VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 VGND VPWR CLK D RESET_B Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_2 VPWR VGND C_N X A B VNB VPB
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.148 ps=1.34 w=0.42 l=0.15
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41o_1 VGND VPWR A3 A4 A2 X B1 A1 VNB VPB
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.184 ps=1.22 w=0.65 l=0.15
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.184 pd=1.22 as=0.161 ps=1.14 w=0.65 l=0.15
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.161 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_4 VPWR VGND X S A1 A0 VNB VPB
X0 a_204_297# A1 a_396_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.16 ps=1.32 w=1 l=0.15
X1 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR S a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_204_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.162 ps=1.33 w=1 l=0.15
X5 a_396_47# A0 a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X6 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.109 ps=0.985 w=0.65 l=0.15
X7 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_490_47# A1 a_396_47# VNB sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.104 ps=0.97 w=0.65 l=0.15
X11 VGND S a_490_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.275 ps=1.5 w=0.65 l=0.15
X12 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_396_47# A0 a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.26 ps=1.45 w=0.65 l=0.15
X14 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VPWR S a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X16 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND S a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 VPWR VGND B D C A X VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_1 VPWR VGND A1 A2 X B1 B2 C1 VNB VPB
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 VPWR VGND A X VNB VPB
X0 a_244_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.217 pd=2.17 as=0.193 ps=1.41 w=0.82 l=0.25
X1 VPWR a_244_47# a_355_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.273 pd=1.61 as=0.217 ps=2.17 w=0.82 l=0.25
X2 X a_355_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.495 pd=2.99 as=0.273 ps=1.61 w=1 l=0.15
X3 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.41 as=0.27 ps=2.54 w=1 l=0.15
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.07 as=0.113 ps=1.38 w=0.42 l=0.15
X5 VGND a_244_47# a_355_47# VNB sky130_fd_pr__nfet_01v8 ad=0.186 pd=1.26 as=0.172 ps=1.83 w=0.65 l=0.25
X6 X a_355_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.83 as=0.186 ps=1.26 w=0.42 l=0.15
X7 a_244_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.123 ps=1.07 w=0.65 l=0.25
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VNB VPB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111o_1 VGND VPWR B1 X D1 A1 A2 C1 VNB VPB
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_2 VGND VPWR X A1 A2 A3 B1 VNB VPB
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.263 ps=2.11 w=0.65 l=0.15
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.175 ps=1.35 w=1 l=0.15
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.405 ps=2.81 w=1 l=0.15
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.213 ps=1.42 w=1 l=0.15
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.114 ps=1 w=0.65 l=0.15
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 VGND VPWR B1_N A1 A2 X VNB VPB
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux4_1 VGND VPWR A1 A0 S0 A3 A2 S1 X VNB VPB
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0852 ps=0.925 w=0.42 l=0.15
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.108 ps=1.36 w=0.42 l=0.15
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.269 pd=2.12 as=0.0921 ps=0.99 w=0.42 l=0.15
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0921 pd=0.99 as=0.109 ps=1.36 w=0.42 l=0.15
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0852 pd=0.925 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0901 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0901 ps=0.995 w=0.42 l=0.15
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.151 ps=1.28 w=0.42 l=0.15
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.151 pd=1.28 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_2 VGND VPWR B C A X VNB VPB
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_1 VGND VPWR B1 B2 A2 A1 X C1 VNB VPB
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.412 pd=1.83 as=0.105 ps=1.21 w=1 l=0.15
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.201 ps=1.92 w=0.65 l=0.15
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0991 ps=0.955 w=0.65 l=0.15
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.412 ps=1.83 w=1 l=0.15
.ends

.subckt Modulator CLK_EXT CLK_PLL CLK_SR Data_SR NMOS1_PS1 NMOS1_PS2 NMOS2_PS1 NMOS2_PS2
+ NMOS_PS3 PMOS1_PS1 PMOS1_PS2 PMOS2_PS1 PMOS2_PS2 PMOS_PS3 RST SIGNAL_OUTPUT VGND
+ VPWR d1[0] d1[1] d1[2] d1[3] d1[4] d1[5] d2[0] d2[1] d2[2] d2[3] d2[4] d2[5]
XFILLER_0_23_247 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1270_ _0626_ _0627_ _0628_ _0512_ VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
X_0985_ VGND VPWR _0442_ _0441_ _0429_ Shift_Register_Inst.data_out\[11\] net23 VGND
+ VPWR sky130_fd_sc_hd__a31o_4
XFILLER_0_1_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0770_ VGND VPWR _0025_ _0280_ _0279_ Signal_Generator_1_90phase_inst.direction _0263_
+ _0281_ VGND VPWR sky130_fd_sc_hd__a32o_1
X_1322_ VPWR VGND Signal_Generator_1_180phase_inst.count\[2\] _0095_ _0009_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_1253_ VGND VPWR _0617_ _0616_ _0513_ _0170_ VGND VPWR sky130_fd_sc_hd__nor3_1
X_1184_ VGND VPWR _0529_ _0558_ _0560_ _0561_ _0559_ VGND VPWR sky130_fd_sc_hd__a22oi_4
XFILLER_0_46_169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0968_ VPWR VGND _0427_ _0424_ _0419_ VGND VPWR sky130_fd_sc_hd__and2_1
X_0899_ VPWR VGND Signal_Generator_2_180phase_inst.count\[2\] _0378_ _0371_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0822_ VPWR VGND _0320_ _0319_ _0310_ _0321_ VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_0_3_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0753_ VGND VPWR Signal_Generator_1_90phase_inst.count\[1\] Signal_Generator_1_90phase_inst.count\[0\]
+ _0268_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0684_ VGND VPWR _0218_ _0216_ _0217_ _0182_ VGND VPWR sky130_fd_sc_hd__mux2_1
X_1305_ VPWR VGND Signal_Generator_1_0phase_inst.direction _0078_ _0006_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_0_36_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1236_ VGND VPWR _0167_ _0603_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1098_ VPWR VGND _0093_ _0515_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1167_ Shift_Register_Inst.data_out\[5\] Shift_Register_Inst.data_out\[6\] _0544_
+ Signal_Generator_1_180phase_inst.count\[3\] VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_19_169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_150 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1021_ VPWR VGND Dead_Time_Generator_inst_1.dt\[2\] _0452_ Dead_Time_Generator_inst_1.dt\[1\]
+ _0455_ _0451_ VGND VPWR sky130_fd_sc_hd__a22o_1
X_0805_ VPWR VGND _0308_ Signal_Generator_1_270phase_inst.count\[0\] Signal_Generator_1_270phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__and2_1
X_0736_ VPWR VGND _0255_ _0254_ _0245_ _0256_ VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_0_24_183 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0667_ VPWR VGND Shift_Register_Inst.shift_state\[0\] _0195_ Shift_Register_Inst.shift_state\[1\]
+ _0205_ VGND VPWR sky130_fd_sc_hd__or3_1
X_1219_ VPWR VGND _0590_ net39 _0587_ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_0_30_120 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xhold30 net55 Signal_Generator_1_180phase_inst.direction VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 net66 Dead_Time_Generator_inst_2.count_dt\[2\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_109 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_125 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1004_ VPWR VGND _0066_ _0449_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_12_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0719_ VPWR VGND _0243_ Signal_Generator_1_0phase_inst.count\[0\] Signal_Generator_1_0phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xoutput20 VGND VPWR net20 PMOS1_PS1 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0984_ VGND VPWR _0441_ _0439_ Shift_Register_Inst.data_out\[12\] clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__and3_4
X_1321_ VPWR VGND Signal_Generator_1_180phase_inst.count\[1\] _0094_ _0008_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1252_ VGND VPWR net37 net29 _0617_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1183_ _0535_ _0541_ _0560_ _0554_ VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_46_137 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0967_ VGND VPWR net22 _0426_ VGND VPWR sky130_fd_sc_hd__buf_1
X_0898_ VPWR VGND Signal_Generator_2_180phase_inst.count\[2\] _0377_ _0374_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_240 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0752_ VGND VPWR _0263_ _0267_ _0027_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0821_ _0320_ Signal_Generator_1_270phase_inst.count\[0\] Signal_Generator_1_270phase_inst.count\[1\]
+ Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[3\]
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_3_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0683_ VGND VPWR _0205_ Shift_Register_Inst.shift_state\[3\] _0187_ _0217_ VGND VPWR
+ sky130_fd_sc_hd__or3b_1
X_1166_ VGND VPWR Shift_Register_Inst.data_out\[5\] Shift_Register_Inst.data_out\[6\]
+ _0543_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1235_ _0601_ _0602_ _0603_ _0561_ VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
X_1304_ Dead_Time_Generator_inst_4.go clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
+ _0157_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_1097_ VPWR VGND _0092_ _0515_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1020_ VGND VPWR _0454_ _0452_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_1.dt\[0\]
+ _0453_ VGND VPWR sky130_fd_sc_hd__o211a_1
X_0735_ _0255_ Signal_Generator_1_0phase_inst.count\[0\] Signal_Generator_1_0phase_inst.count\[1\]
+ Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[3\]
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
X_0804_ _0307_ Signal_Generator_1_270phase_inst.count\[5\] Signal_Generator_1_270phase_inst.count\[4\]
+ _0305_ _0306_ VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
X_0666_ VGND VPWR _0149_ _0204_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1149_ VGND VPWR Shift_Register_Inst.data_out\[16\] _0526_ net7 VGND VPWR sky130_fd_sc_hd__or2b_1
XFILLER_0_27_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1218_ VGND VPWR _0584_ _0586_ _0588_ _0589_ VGND VPWR sky130_fd_sc_hd__o21a_1
Xhold42 net67 Shift_Register_Inst.data_out\[17\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 net45 Dead_Time_Generator_inst_3.count_dt\[3\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 net56 Dead_Time_Generator_inst_1.count_dt\[0\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1003_ VPWR VGND _0449_ _0446_ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_12_110 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0718_ _0242_ Signal_Generator_1_0phase_inst.count\[5\] Signal_Generator_1_0phase_inst.count\[4\]
+ _0240_ _0241_ VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
X_0649_ VPWR VGND _0193_ _0192_ _0189_ VGND VPWR sky130_fd_sc_hd__and2_1
Xoutput21 VGND VPWR net21 PMOS1_PS2 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_202 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0983_ VGND VPWR _0440_ _0432_ _0438_ net18 _0439_ VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_0_22_271 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_6 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1320_ VPWR VGND Signal_Generator_1_180phase_inst.count\[0\] _0093_ _0007_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1182_ VPWR VGND _0540_ _0539_ _0559_ _0557_ _0528_ VGND VPWR sky130_fd_sc_hd__a211oi_2
X_1251_ VPWR VGND _0616_ _0615_ Dead_Time_Generator_inst_3.count_dt\[0\] VGND VPWR
+ sky130_fd_sc_hd__and2_1
XFILLER_0_24_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0897_ VPWR VGND _0375_ _0041_ _0376_ _0036_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0966_ VGND VPWR _0417_ _0424_ _0416_ _0426_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_4_51 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_216 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0751_ VGND VPWR _0267_ Signal_Generator_1_90phase_inst.count\[4\] net53 _0266_ VGND
+ VPWR sky130_fd_sc_hd__and3_1
X_0820_ VPWR VGND _0319_ _0309_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_10_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0682_ VGND VPWR Shift_Register_Inst.data_out\[8\] _0216_ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_1303_ VGND VPWR clknet_1_1__leaf_CLK_SR _0156_ _0077_ Shift_Register_Inst.shift_state\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1096_ VPWR VGND _0091_ _0515_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1165_ VGND VPWR Shift_Register_Inst.data_out\[13\] _0542_ net6 VGND VPWR sky130_fd_sc_hd__or2b_1
X_1234_ _0602_ _0594_ Dead_Time_Generator_inst_2.count_dt\[1\] Dead_Time_Generator_inst_2.count_dt\[2\]
+ Dead_Time_Generator_inst_2.count_dt\[3\] VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
X_0949_ VGND VPWR _0414_ net5 _0228_ Dead_Time_Generator_inst_4.go VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_33_130 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0734_ VPWR VGND _0254_ _0244_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0803_ VPWR VGND _0306_ Signal_Generator_1_270phase_inst.direction VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_24_141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0665_ VGND VPWR _0204_ Dead_Time_Generator_inst_1.dt\[3\] _0203_ _0182_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
X_1148_ VGND VPWR _0525_ _0519_ _0524_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1217_ VGND VPWR _0587_ Dead_Time_Generator_inst_1.dt\[2\] _0585_ Dead_Time_Generator_inst_1.dt\[3\]
+ _0588_ VGND VPWR sky130_fd_sc_hd__o22a_1
X_1079_ VPWR VGND _0513_ _0512_ VGND VPWR sky130_fd_sc_hd__buf_2
Xhold21 net46 Signal_Generator_2_90phase_inst.count\[0\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 net68 Signal_Generator_2_180phase_inst.direction VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 net35 Signal_Generator_1_270phase_inst.count\[0\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 net57 Shift_Register_Inst.shift_state\[1\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_244 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1002_ VPWR VGND _0065_ _0448_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0717_ VPWR VGND _0241_ Signal_Generator_1_0phase_inst.direction VGND VPWR sky130_fd_sc_hd__inv_2
X_0648_ VGND VPWR _0192_ _0187_ _0188_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_35_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput22 VGND VPWR net22 PMOS2_PS1 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0982_ VPWR VGND _0439_ Shift_Register_Inst.data_out\[11\] VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_13_250 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1181_ VPWR VGND _0556_ _0555_ _0557_ _0558_ VGND VPWR sky130_fd_sc_hd__a21o_1
X_1250_ _0615_ _0611_ _0612_ _0613_ net28 VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_24_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0896_ VPWR VGND _0375_ _0370_ net51 _0376_ VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_269 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0965_ VGND VPWR net15 _0425_ VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_4_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1379_ Dead_Time_Generator_inst_4.count_dt\[0\] clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
+ _0176_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0750_ VGND VPWR _0266_ Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[3\]
+ _0265_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0681_ VGND VPWR _0145_ _0215_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1302_ VGND VPWR clknet_1_1__leaf_CLK_SR _0155_ _0076_ Shift_Register_Inst.shift_state\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1233_ VGND VPWR _0601_ Dead_Time_Generator_inst_2.count_dt\[2\] Dead_Time_Generator_inst_2.count_dt\[3\]
+ _0597_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1095_ VPWR VGND _0090_ _0515_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1164_ VPWR VGND _0541_ _0228_ _0530_ _0534_ _0540_ _0539_ VGND VPWR sky130_fd_sc_hd__o32a_1
XFILLER_0_27_172 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0948_ VGND VPWR Shift_Register_Inst.data_out\[16\] Shift_Register_Inst.data_out\[17\]
+ Shift_Register_Inst.data_out\[15\] _0413_ VGND VPWR sky130_fd_sc_hd__or3b_1
X_0879_ VPWR VGND _0363_ _0349_ _0360_ _0052_ net52 VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_0_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_142 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0802_ VPWR VGND Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[0\]
+ Signal_Generator_1_270phase_inst.count\[1\] Signal_Generator_1_270phase_inst.count\[3\]
+ _0305_ VGND VPWR sky130_fd_sc_hd__or4_2
X_0733_ VGND VPWR _0240_ _0253_ _0252_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_0664_ VGND VPWR _0187_ _0188_ _0186_ _0203_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_21_98 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1216_ VPWR VGND _0587_ Dead_Time_Generator_inst_2.count_dt\[3\] VGND VPWR sky130_fd_sc_hd__inv_2
X_1078_ _0512_ _0477_ _0494_ _0507_ _0511_ VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
X_1147_ VGND VPWR _0523_ _0520_ Signal_Generator_1_0phase_inst.count\[5\] _0521_ _0524_
+ VGND VPWR sky130_fd_sc_hd__o22a_1
Xhold22 net47 Signal_Generator_2_180phase_inst.count\[0\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 net36 Dead_Time_Generator_inst_1.count_dt\[4\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 net69 Signal_Generator_2_0phase_inst.direction VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 net58 Signal_Generator_1_0phase_inst.direction VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_1001_ VPWR VGND _0064_ _0448_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_16_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0716_ VPWR VGND Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[0\]
+ Signal_Generator_1_0phase_inst.count\[1\] Signal_Generator_1_0phase_inst.count\[3\]
+ _0240_ VGND VPWR sky130_fd_sc_hd__or4_2
X_0647_ VGND VPWR _0190_ _0155_ _0191_ VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_0_35_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput23 VGND VPWR net23 PMOS2_PS2 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_194 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_218 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0981_ VPWR VGND _0430_ net21 _0437_ _0438_ VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_0_1_145 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_189 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1180_ VGND VPWR _0527_ _0525_ _0557_ _0526_ VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0964_ VPWR VGND _0425_ _0424_ _0414_ VGND VPWR sky130_fd_sc_hd__and2_1
X_0895_ VGND VPWR _0375_ _0374_ _0371_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_10_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1378_ Dead_Time_Generator_inst_2.go clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
+ _0175_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0680_ VGND VPWR _0215_ _0214_ _0190_ _0182_ VGND VPWR sky130_fd_sc_hd__mux2_1
X_1301_ VGND VPWR clknet_1_1__leaf_CLK_SR _0154_ _0075_ Shift_Register_Inst.shift_state\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1232_ VGND VPWR _0581_ _0600_ _0166_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1094_ VPWR VGND _0089_ _0515_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1163_ VGND VPWR _0228_ _0540_ net3 VGND VPWR sky130_fd_sc_hd__or2b_1
X_0947_ VPWR VGND net24 _0412_ VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_27_162 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0878_ VPWR VGND _0362_ _0361_ _0352_ _0363_ VGND VPWR sky130_fd_sc_hd__a21o_1
X_0801_ _0012_ _0287_ Signal_Generator_1_180phase_inst.direction Signal_Generator_1_180phase_inst.count\[4\]
+ _0304_ VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_24_132 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0732_ Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[1\]
+ Signal_Generator_1_0phase_inst.count\[0\] _0252_ Signal_Generator_1_0phase_inst.count\[3\]
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31ai_1
X_0663_ VGND VPWR _0150_ _0202_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1146_ _0523_ Signal_Generator_1_270phase_inst.count\[5\] _0211_ _0208_ _0522_ VGND
+ VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
X_1215_ VPWR VGND Dead_Time_Generator_inst_1.dt\[2\] _0582_ Dead_Time_Generator_inst_1.dt\[1\]
+ _0586_ _0585_ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_1_76 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1077_ VGND VPWR _0475_ _0477_ _0510_ _0511_ _0476_ VGND VPWR sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_15_165 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_121 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xhold34 net59 Signal_Generator_2_0phase_inst.direction VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 net37 Dead_Time_Generator_inst_3.count_dt\[0\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 net48 Shift_Register_Inst.shift_state\[4\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_1000_ VPWR VGND _0063_ _0448_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_16_99 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0715_ VGND VPWR _0135_ _0239_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0646_ VGND VPWR _0186_ _0191_ _0189_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_1129_ VPWR VGND _0121_ _0518_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_35_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput24 VGND VPWR net24 PMOS_PS3 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_75 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0980_ VGND VPWR _0437_ Shift_Register_Inst.data_out\[10\] Shift_Register_Inst.data_out\[9\]
+ net16 VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_1_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_0__f_Dead_Time_Generator_inst_1.clk VGND VPWR clknet_0_Dead_Time_Generator_inst_1.clk
+ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_0894_ VGND VPWR Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_180phase_inst.count\[1\]
+ _0374_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_6_205 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0963_ Shift_Register_Inst.data_out\[16\] Shift_Register_Inst.data_out\[17\] _0424_
+ Shift_Register_Inst.data_out\[15\] VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_4_43 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1377_ Dead_Time_Generator_inst_3.count_dt\[4\] clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
+ _0174_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_1162_ VPWR VGND _0539_ _0536_ _0537_ _0538_ Signal_Generator_1_0phase_inst.count\[0\]
+ _0520_ VGND VPWR sky130_fd_sc_hd__o32a_1
X_1231_ VGND VPWR _0597_ _0600_ net66 VGND VPWR sky130_fd_sc_hd__xnor2_1
X_1300_ VGND VPWR clknet_1_0__leaf_CLK_SR _0153_ _0074_ Shift_Register_Inst.shift_state\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1093_ VPWR VGND _0088_ _0515_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0877_ _0362_ Signal_Generator_2_90phase_inst.count\[2\] Signal_Generator_2_90phase_inst.count\[1\]
+ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[3\]
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
X_0946_ VGND VPWR net7 _0412_ Shift_Register_Inst.data_out\[16\] VGND VPWR sky130_fd_sc_hd__or2b_1
XFILLER_0_27_152 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0731_ VPWR VGND _0251_ _0242_ _0249_ _0002_ Signal_Generator_1_0phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__a22o_1
X_0800_ _0304_ Signal_Generator_1_180phase_inst.count\[4\] Signal_Generator_1_180phase_inst.direction
+ _0283_ Signal_Generator_1_180phase_inst.count\[5\] VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
X_0662_ VGND VPWR _0202_ Dead_Time_Generator_inst_1.dt\[2\] _0201_ _0182_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1145_ _0211_ Signal_Generator_1_90phase_inst.count\[5\] _0522_ _0208_ VGND VPWR
+ VGND VPWR sky130_fd_sc_hd__and3b_1
X_1214_ VPWR VGND _0585_ Dead_Time_Generator_inst_2.count_dt\[2\] VGND VPWR sky130_fd_sc_hd__inv_2
X_1076_ VGND VPWR _0509_ _0492_ _0508_ _0494_ _0510_ VGND VPWR sky130_fd_sc_hd__o22a_1
X_0929_ VPWR VGND _0400_ _0391_ _0398_ _0044_ Signal_Generator_2_270phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_15_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold13 net38 _0170_ VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 net49 Dead_Time_Generator_inst_1.count_dt\[1\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 net60 Shift_Register_Inst.shift_state\[0\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_158 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_203 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0645_ VGND VPWR _0190_ _0186_ _0189_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0714_ VGND VPWR _0239_ net1 _0238_ net67 VGND VPWR sky130_fd_sc_hd__mux2_1
X_1128_ VPWR VGND _0120_ _0518_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1059_ VPWR VGND _0490_ _0489_ _0485_ _0493_ VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_174 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput25 VGND VPWR net25 SIGNAL_OUTPUT VGND VPWR sky130_fd_sc_hd__buf_8
XPHY_0 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_242 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_220 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0893_ VPWR VGND _0035_ net47 VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_6_217 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0962_ VPWR VGND net21 _0423_ VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
X_1376_ Dead_Time_Generator_inst_3.count_dt\[3\] clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
+ _0173_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_14 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1161_ VGND VPWR _0208_ _0007_ _0538_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1092_ VPWR VGND _0087_ _0515_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1230_ VGND VPWR _0165_ _0599_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0876_ VPWR VGND _0361_ _0351_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_42_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0945_ VGND VPWR _0411_ net19 VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_1359_ VGND VPWR clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0046_ _0132_ Signal_Generator_2_270phase_inst.count\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_153 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0730_ VGND VPWR _0251_ _0245_ _0250_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0661_ VPWR VGND _0187_ _0200_ Shift_Register_Inst.shift_state\[3\] _0201_ VGND VPWR
+ sky130_fd_sc_hd__or3_1
X_1213_ VGND VPWR _0584_ _0582_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_1.dt\[0\]
+ _0583_ VGND VPWR sky130_fd_sc_hd__o211a_1
X_1075_ VPWR VGND _0504_ _0503_ _0506_ _0509_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_1144_ VPWR VGND _0300_ _0211_ _0208_ _0521_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0859_ VPWR VGND _0348_ Signal_Generator_2_90phase_inst.direction VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_30_137 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0928_ VGND VPWR _0400_ _0394_ _0399_ VGND VPWR sky130_fd_sc_hd__or2_1
Xhold36 net61 Signal_Generator_1_270phase_inst.direction VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 net50 Dead_Time_Generator_inst_3.count_dt\[1\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 net39 Dead_Time_Generator_inst_1.dt\[3\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_215 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_137 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0644_ VGND VPWR _0187_ _0189_ _0188_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_0713_ VGND VPWR _0238_ Shift_Register_Inst.shift_state\[0\] Shift_Register_Inst.shift_state\[4\]
+ _0237_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_32_6 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1127_ VPWR VGND _0119_ _0518_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1058_ VPWR VGND _0483_ _0482_ _0478_ _0492_ VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_186 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput15 VGND VPWR net15 NMOS1_PS1 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_34 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_262 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0961_ VGND VPWR _0423_ _0413_ _0422_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0892_ VGND VPWR _0370_ _0373_ _0041_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_6_229 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_45 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1375_ Dead_Time_Generator_inst_3.count_dt\[2\] clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
+ _0172_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_132 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_37 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1160_ VPWR VGND _0021_ _0208_ _0211_ _0537_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_1091_ VPWR VGND _0086_ _0515_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_35_67 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0944_ VPWR VGND _0411_ net8 Shift_Register_Inst.data_out\[16\] VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_0_2_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0875_ VGND VPWR _0347_ _0360_ _0359_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_1358_ VGND VPWR clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0045_ _0131_ Signal_Generator_2_270phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1289_ VGND VPWR clknet_1_1__leaf_CLK_SR _0142_ _0063_ Shift_Register_Inst.data_out\[10\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_176 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0660_ VPWR VGND Shift_Register_Inst.shift_state\[1\] _0200_ Shift_Register_Inst.shift_state\[4\]
+ Shift_Register_Inst.shift_state\[0\] VGND VPWR sky130_fd_sc_hd__or3b_2
XFILLER_0_46_66 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1212_ VPWR VGND _0583_ Dead_Time_Generator_inst_2.count_dt\[0\] VGND VPWR sky130_fd_sc_hd__inv_2
X_1074_ VGND VPWR _0484_ _0491_ _0508_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1143_ VGND VPWR _0520_ Shift_Register_Inst.data_out\[5\] Shift_Register_Inst.data_out\[6\]
+ VGND VPWR sky130_fd_sc_hd__or2_1
X_0927_ VPWR VGND Signal_Generator_2_270phase_inst.count\[2\] _0399_ _0392_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_157 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0858_ VPWR VGND Signal_Generator_2_90phase_inst.count\[1\] Signal_Generator_2_90phase_inst.count\[2\]
+ Signal_Generator_2_90phase_inst.count\[3\] Signal_Generator_2_90phase_inst.count\[0\]
+ _0347_ VGND VPWR sky130_fd_sc_hd__or4_2
X_0789_ Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[1\]
+ Signal_Generator_1_180phase_inst.count\[0\] _0295_ Signal_Generator_1_180phase_inst.count\[3\]
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31ai_1
Xhold26 VGND VPWR net51 Signal_Generator_2_180phase_inst.direction VGND VPWR sky130_fd_sc_hd__buf_1
Xhold15 net40 Dead_Time_Generator_inst_1.count_dt\[3\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 net62 Dead_Time_Generator_inst_3.count_dt\[2\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_260 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_260 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0643_ Shift_Register_Inst.shift_state\[4\] Shift_Register_Inst.shift_state\[1\]
+ _0188_ Shift_Register_Inst.shift_state\[0\] VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
X_0712_ VPWR VGND _0237_ _0183_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1126_ VPWR VGND _0118_ _0518_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1057_ VGND VPWR _0491_ _0489_ _0485_ _0490_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_7_154 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput16 VGND VPWR net16 NMOS1_PS2 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_219 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_45 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_208 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_274 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1109_ VPWR VGND _0103_ _0516_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_23_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_274 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_67 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0960_ VGND VPWR _0422_ net6 _0228_ _0421_ VGND VPWR sky130_fd_sc_hd__mux2_1
X_0891_ VGND VPWR _0373_ Signal_Generator_2_180phase_inst.count\[4\] Signal_Generator_2_180phase_inst.count\[5\]
+ _0372_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_40_68 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1374_ Dead_Time_Generator_inst_3.count_dt\[1\] clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
+ _0171_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_144 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_122 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1090_ VPWR VGND _0515_ _0446_ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_35_79 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0874_ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[1\]
+ Signal_Generator_2_90phase_inst.count\[2\] _0359_ Signal_Generator_2_90phase_inst.count\[3\]
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31ai_1
X_0943_ VPWR VGND Dead_Time_Generator_inst_1.clk _0410_ VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_0_2_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1288_ VGND VPWR clknet_1_1__leaf_CLK_SR _0141_ _0062_ Shift_Register_Inst.data_out\[11\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1357_ VGND VPWR clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0044_ _0130_ Signal_Generator_2_270phase_inst.count\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_188 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_78 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1142_ VGND VPWR Shift_Register_Inst.data_out\[16\] _0519_ net8 VGND VPWR sky130_fd_sc_hd__or2b_1
X_1211_ VPWR VGND _0582_ Dead_Time_Generator_inst_2.count_dt\[1\] VGND VPWR sky130_fd_sc_hd__inv_2
X_1073_ VGND VPWR _0507_ _0496_ _0505_ _0495_ _0506_ VGND VPWR sky130_fd_sc_hd__a211o_1
X_0857_ _0033_ _0330_ Signal_Generator_2_0phase_inst.direction net65 _0346_ VGND VPWR
+ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0926_ VPWR VGND Signal_Generator_2_270phase_inst.count\[2\] _0398_ _0395_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold27 VGND VPWR net52 Signal_Generator_2_90phase_inst.direction VGND VPWR sky130_fd_sc_hd__buf_1
X_0788_ VPWR VGND _0294_ _0285_ _0292_ _0009_ net55 VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold16 net41 _0580_ VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 net63 Dead_Time_Generator_inst_1.count_dt\[2\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_69 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0711_ VGND VPWR _0136_ _0236_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_1__f_Dead_Time_Generator_inst_1.clk VGND VPWR clknet_0_Dead_Time_Generator_inst_1.clk
+ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_0642_ VGND VPWR Shift_Register_Inst.shift_state\[1\] Shift_Register_Inst.shift_state\[0\]
+ _0187_ _0156_ net48 _0186_ VGND VPWR sky130_fd_sc_hd__a41o_1
X_1125_ VPWR VGND _0117_ _0518_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1056_ VGND VPWR _0490_ Signal_Generator_2_0phase_inst.count\[2\] _0467_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_0909_ VGND VPWR _0386_ Signal_Generator_2_180phase_inst.count\[4\] _0372_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
Xoutput17 VGND VPWR net17 NMOS2_PS1 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_223 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1039_ VGND VPWR _0473_ _0216_ _0214_ Signal_Generator_2_270phase_inst.count\[5\]
+ VGND VPWR sky130_fd_sc_hd__and3_1
X_1108_ VPWR VGND _0102_ _0516_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_16_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_220 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_57 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0890_ VGND VPWR _0372_ Signal_Generator_2_180phase_inst.count\[2\] Signal_Generator_2_180phase_inst.count\[3\]
+ _0371_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1373_ Dead_Time_Generator_inst_3.count_dt\[0\] clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
+ net38 VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_156 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_134 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0873_ VPWR VGND _0358_ _0349_ _0356_ _0051_ net52 VGND VPWR sky130_fd_sc_hd__a22o_1
X_0942_ VPWR VGND _0410_ Shift_Register_Inst.data_out\[14\] CLK_EXT CLK_PLL VGND VPWR
+ sky130_fd_sc_hd__mux2_4
XFILLER_0_2_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1287_ VGND VPWR clknet_1_1__leaf_CLK_SR _0140_ _0061_ Shift_Register_Inst.data_out\[12\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1356_ VGND VPWR clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0043_ _0129_ Signal_Generator_2_270phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1072_ VGND VPWR _0506_ _0497_ _0502_ _0501_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_46_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_35 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1210_ VPWR VGND _0134_ _0447_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1141_ VPWR VGND _0133_ _0447_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0856_ _0346_ Signal_Generator_2_0phase_inst.count\[4\] Signal_Generator_2_0phase_inst.direction
+ _0326_ Signal_Generator_2_0phase_inst.count\[5\] VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
X_0787_ VGND VPWR _0294_ _0288_ _0293_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_30_129 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0925_ VPWR VGND _0396_ _0048_ _0397_ _0043_ VGND VPWR sky130_fd_sc_hd__a21oi_1
Xhold28 net53 Signal_Generator_1_90phase_inst.count\[5\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold17 net42 Signal_Generator_1_0phase_inst.count\[0\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 net64 Shift_Register_Inst.data_out\[15\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_1339_ VGND VPWR clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0033_ _0112_ Signal_Generator_2_0phase_inst.count\[5\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_0641_ VGND VPWR Shift_Register_Inst.shift_state\[2\] _0187_ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_0710_ VGND VPWR _0236_ Shift_Register_Inst.data_out\[16\] _0235_ net1 VGND VPWR
+ sky130_fd_sc_hd__mux2_1
X_1124_ VPWR VGND _0116_ _0518_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1055_ VPWR VGND _0486_ _0488_ _0487_ _0471_ _0489_ VGND VPWR sky130_fd_sc_hd__or4_1
Xoutput18 VGND VPWR net18 NMOS2_PS2 VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_0839_ VGND VPWR _0333_ _0332_ _0329_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0908_ VGND VPWR Signal_Generator_2_180phase_inst.count\[5\] Signal_Generator_2_180phase_inst.count\[4\]
+ _0382_ _0385_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_19_240 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1038_ VPWR VGND Signal_Generator_2_90phase_inst.count\[5\] _0463_ _0472_ _0464_
+ Signal_Generator_2_180phase_inst.count\[5\] _0471_ VGND VPWR sky130_fd_sc_hd__a221o_1
X_1107_ VPWR VGND _0101_ _0516_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_17_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_202 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_216 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_37 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1372_ Dead_Time_Generator_inst_1.go clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
+ _0169_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0941_ _0047_ _0393_ Signal_Generator_2_270phase_inst.direction Signal_Generator_2_270phase_inst.count\[4\]
+ _0409_ VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
X_0872_ VGND VPWR _0358_ _0352_ _0357_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1355_ VGND VPWR clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0042_ _0128_ Signal_Generator_2_270phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1286_ VGND VPWR clknet_1_0__leaf_CLK_SR _0139_ _0060_ Shift_Register_Inst.data_out\[13\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_91 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1071_ VGND VPWR _0503_ _0505_ _0504_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_1140_ VPWR VGND _0132_ _0447_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_46_47 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0924_ VPWR VGND _0396_ _0391_ Signal_Generator_2_270phase_inst.direction _0397_
+ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0855_ VGND VPWR _0032_ _0344_ _0343_ Signal_Generator_2_0phase_inst.direction _0328_
+ _0345_ VGND VPWR sky130_fd_sc_hd__a32o_1
X_0786_ VPWR VGND Signal_Generator_1_180phase_inst.count\[2\] _0293_ _0286_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_108 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1338_ VGND VPWR clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0032_ _0111_ Signal_Generator_2_0phase_inst.count\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
Xhold18 net43 Signal_Generator_1_90phase_inst.count\[0\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 VPWR VGND Signal_Generator_1_90phase_inst.direction net54 VGND VPWR sky130_fd_sc_hd__clkdlybuf4s25_1
X_1269_ VGND VPWR _0627_ Dead_Time_Generator_inst_4.count_dt\[1\] _0623_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
XFILLER_0_21_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_160 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_49 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0640_ VPWR VGND _0186_ Shift_Register_Inst.shift_state\[3\] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_20_141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1123_ VPWR VGND _0518_ _0446_ VGND VPWR sky130_fd_sc_hd__buf_4
X_1054_ VGND VPWR _0488_ Shift_Register_Inst.data_out\[8\] Shift_Register_Inst.data_out\[7\]
+ Signal_Generator_2_270phase_inst.count\[2\] VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_7_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0907_ VPWR VGND _0384_ _0370_ _0381_ _0038_ net51 VGND VPWR sky130_fd_sc_hd__a22o_1
X_0838_ VGND VPWR Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[1\]
+ _0332_ VGND VPWR sky130_fd_sc_hd__nor2_1
Xoutput19 VGND VPWR net19 NMOS_PS3 VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_0769_ VGND VPWR _0261_ _0281_ Signal_Generator_1_90phase_inst.count\[4\] VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1106_ VPWR VGND _0100_ _0516_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1037_ VGND VPWR Shift_Register_Inst.data_out\[7\] Shift_Register_Inst.data_out\[8\]
+ _0471_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_17_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_266 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_269 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_155 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_228 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1371_ Dead_Time_Generator_inst_2.count_dt\[4\] clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk
+ _0168_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0940_ _0409_ Signal_Generator_2_270phase_inst.count\[4\] Signal_Generator_2_270phase_inst.direction
+ _0389_ Signal_Generator_2_270phase_inst.count\[5\] VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
X_0871_ VPWR VGND Signal_Generator_2_90phase_inst.count\[2\] _0357_ _0350_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1285_ VGND VPWR clknet_1_0__leaf_CLK_SR _0138_ _0059_ Shift_Register_Inst.data_out\[14\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1354_ VGND VPWR clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0048_ _0127_ Signal_Generator_2_270phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_114 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1070_ VGND VPWR _0504_ _0495_ _0496_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0854_ VGND VPWR _0326_ _0345_ Signal_Generator_2_0phase_inst.count\[4\] VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0923_ VGND VPWR _0396_ _0395_ _0392_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0785_ VPWR VGND Signal_Generator_1_180phase_inst.count\[2\] _0292_ _0289_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_172 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_150 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1337_ VGND VPWR clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0031_ _0110_ Signal_Generator_2_0phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xhold19 net44 Signal_Generator_1_180phase_inst.count\[0\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_1268_ VGND VPWR _0626_ Dead_Time_Generator_inst_4.count_dt\[0\] Dead_Time_Generator_inst_4.count_dt\[1\]
+ _0461_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1199_ VGND VPWR _0575_ _0574_ _0561_ _0158_ VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_0_14_172 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1122_ VPWR VGND _0115_ _0517_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1053_ Shift_Register_Inst.data_out\[8\] Signal_Generator_2_90phase_inst.count\[2\]
+ _0487_ Shift_Register_Inst.data_out\[7\] VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
X_0837_ VPWR VGND _0028_ net34 VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_7_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0906_ VPWR VGND _0383_ _0382_ _0373_ _0384_ VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_0_28_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_94 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0768_ VGND VPWR _0280_ Signal_Generator_1_90phase_inst.count\[4\] _0266_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_0699_ VPWR VGND _0228_ Shift_Register_Inst.data_out\[13\] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_34_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1105_ VPWR VGND _0099_ _0516_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_16_6 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1036_ VPWR VGND _0470_ net14 VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_3_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1019_ VPWR VGND _0453_ Dead_Time_Generator_inst_4.count_dt\[0\] VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_8_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1370_ Dead_Time_Generator_inst_2.count_dt\[3\] clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk
+ _0167_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0870_ VPWR VGND Signal_Generator_2_90phase_inst.count\[2\] _0356_ _0353_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
Xclkbuf_3_2__f_Dead_Time_Generator_inst_1.clk VGND VPWR clknet_0_Dead_Time_Generator_inst_1.clk
+ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_1353_ VPWR VGND Signal_Generator_2_180phase_inst.count\[5\] _0126_ _0040_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1284_ VGND VPWR clknet_1_0__leaf_CLK_SR _0137_ _0058_ Shift_Register_Inst.data_out\[15\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_140 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0999_ VPWR VGND _0062_ _0448_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_33_118 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0853_ VGND VPWR _0344_ Signal_Generator_2_0phase_inst.count\[4\] _0330_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_0922_ VGND VPWR Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[1\]
+ _0395_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0784_ VPWR VGND _0290_ _0013_ _0291_ _0008_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_1336_ VGND VPWR clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0030_ _0109_ Signal_Generator_2_0phase_inst.count\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
Xinput1 VPWR VGND net1 Data_SR VGND VPWR sky130_fd_sc_hd__buf_2
X_1198_ VGND VPWR net56 _0573_ _0575_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1267_ VGND VPWR _0176_ _0625_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_221 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_184 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_154 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1121_ VPWR VGND _0114_ _0517_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1052_ Shift_Register_Inst.data_out\[7\] Shift_Register_Inst.data_out\[8\] _0486_
+ Signal_Generator_2_180phase_inst.count\[2\] VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_7_137 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0836_ VGND VPWR _0328_ _0331_ _0034_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0905_ _0383_ Signal_Generator_2_180phase_inst.count\[2\] Signal_Generator_2_180phase_inst.count\[1\]
+ Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_180phase_inst.count\[3\]
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
X_0767_ VGND VPWR Signal_Generator_1_90phase_inst.count\[5\] Signal_Generator_1_90phase_inst.count\[4\]
+ _0276_ _0279_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_44_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0698_ VGND VPWR _0140_ _0227_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1319_ VPWR VGND Signal_Generator_1_180phase_inst.direction _0092_ _0013_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
XPHY_7 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1035_ VGND VPWR _0462_ _0468_ _0469_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1104_ VPWR VGND _0098_ _0516_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_17_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0819_ VGND VPWR _0305_ _0318_ _0317_ VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_0_31_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1018_ VPWR VGND _0452_ Dead_Time_Generator_inst_4.count_dt\[1\] VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_8_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_116 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1352_ VPWR VGND Signal_Generator_2_180phase_inst.count\[4\] _0125_ _0039_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_1283_ VGND VPWR clknet_1_0__leaf_CLK_SR _0136_ _0057_ Shift_Register_Inst.data_out\[16\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0998_ VPWR VGND _0061_ _0448_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_24_119 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0921_ VPWR VGND _0042_ net32 VGND VPWR sky130_fd_sc_hd__inv_2
X_0852_ VGND VPWR Signal_Generator_2_0phase_inst.count\[5\] Signal_Generator_2_0phase_inst.count\[4\]
+ _0340_ _0343_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_11_86 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0783_ VPWR VGND _0290_ _0285_ net55 _0291_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_1335_ VGND VPWR clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0029_ _0108_ Signal_Generator_2_0phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput2 VGND VPWR net2 RST VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_72 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1197_ VPWR VGND _0574_ _0573_ Dead_Time_Generator_inst_1.count_dt\[0\] VGND VPWR
+ sky130_fd_sc_hd__and2_1
X_1266_ _0623_ _0624_ _0625_ _0513_ VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_20_166 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1120_ VPWR VGND _0113_ _0517_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1051_ VPWR VGND _0485_ net11 VGND VPWR sky130_fd_sc_hd__inv_2
X_0904_ VPWR VGND _0382_ _0372_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_43_203 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0835_ VGND VPWR _0331_ Signal_Generator_2_0phase_inst.count\[4\] Signal_Generator_2_0phase_inst.count\[5\]
+ _0330_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0766_ VPWR VGND _0278_ _0263_ _0275_ _0024_ net54 VGND VPWR sky130_fd_sc_hd__a22o_1
X_0697_ VGND VPWR _0227_ Shift_Register_Inst.data_out\[12\] _0226_ net1 VGND VPWR
+ sky130_fd_sc_hd__mux2_1
X_1318_ VGND VPWR clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0026_ _0091_ Signal_Generator_1_90phase_inst.count\[5\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1249_ VGND VPWR net27 _0614_ Dead_Time_Generator_inst_3.count_dt\[4\] VGND VPWR
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_6_182 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1034_ VGND VPWR _0468_ _0466_ _0467_ Signal_Generator_2_0phase_inst.count\[4\] VGND
+ VPWR sky130_fd_sc_hd__mux2_1
X_1103_ VPWR VGND _0097_ _0516_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_31_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0749_ VGND VPWR _0264_ _0021_ _0265_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0818_ Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[1\]
+ Signal_Generator_1_270phase_inst.count\[0\] _0317_ Signal_Generator_1_270phase_inst.count\[3\]
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31ai_1
XFILLER_0_38_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1017_ VPWR VGND _0451_ Dead_Time_Generator_inst_4.count_dt\[2\] VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_39_125 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_150 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_180 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1351_ VPWR VGND Signal_Generator_2_180phase_inst.count\[3\] _0124_ _0038_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_0_25_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1282_ VGND VPWR clknet_1_0__leaf_CLK_SR _0135_ _0056_ Shift_Register_Inst.data_out\[17\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0997_ VPWR VGND _0060_ _0448_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_17_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0920_ VGND VPWR _0391_ _0394_ _0048_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0851_ VPWR VGND _0342_ _0328_ _0339_ _0031_ Signal_Generator_2_0phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_11_98 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0782_ VGND VPWR _0290_ _0289_ _0286_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1334_ VGND VPWR clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0028_ _0107_ Signal_Generator_2_0phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1265_ VGND VPWR _0624_ Dead_Time_Generator_inst_4.count_dt\[0\] _0461_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_1196_ _0573_ _0569_ _0570_ _0571_ _0572_ VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
Xinput3 VGND VPWR net3 d1[0] VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_14_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1050_ VGND VPWR _0484_ _0482_ _0478_ _0483_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0834_ VGND VPWR _0330_ Signal_Generator_2_0phase_inst.count\[2\] Signal_Generator_2_0phase_inst.count\[3\]
+ _0329_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_7_106 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0903_ VGND VPWR _0368_ _0381_ _0380_ VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_0_43_215 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0765_ VPWR VGND _0277_ _0276_ _0267_ _0278_ VGND VPWR sky130_fd_sc_hd__a21o_1
X_0696_ VGND VPWR _0226_ _0225_ _0205_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1317_ VPWR VGND Signal_Generator_1_90phase_inst.count\[4\] _0090_ _0025_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_1248_ _0613_ Dead_Time_Generator_inst_3.count_dt\[4\] net27 VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__and2b_1
X_1179_ VGND VPWR _0551_ _0556_ _0552_ VGND VPWR sky130_fd_sc_hd__nand2_1
XPHY_9 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_207 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1102_ VPWR VGND _0096_ _0516_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1033_ VGND VPWR _0467_ _0214_ _0216_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0817_ VPWR VGND _0316_ _0307_ _0314_ _0016_ Signal_Generator_1_270phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_24_270 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0679_ VGND VPWR Shift_Register_Inst.data_out\[7\] _0214_ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_0748_ VPWR VGND _0021_ net43 VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_0_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1016_ VPWR VGND _0077_ _0450_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_5_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_107 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1350_ VPWR VGND Signal_Generator_2_180phase_inst.count\[2\] _0123_ _0037_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_1281_ VGND VPWR _0513_ net29 _0181_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0996_ VPWR VGND _0059_ _0448_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_1_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0850_ VPWR VGND _0341_ _0340_ _0331_ _0342_ VGND VPWR sky130_fd_sc_hd__a21o_1
X_0781_ VGND VPWR Signal_Generator_1_180phase_inst.count\[1\] Signal_Generator_1_180phase_inst.count\[0\]
+ _0289_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1333_ VPWR VGND Signal_Generator_2_0phase_inst.direction _0106_ _0034_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
Xinput4 VGND VPWR net4 d1[1] VGND VPWR sky130_fd_sc_hd__buf_1
X_1264_ VPWR VGND _0623_ _0461_ Dead_Time_Generator_inst_4.count_dt\[0\] VGND VPWR
+ sky130_fd_sc_hd__and2_1
X_1195_ VGND VPWR net27 _0572_ Dead_Time_Generator_inst_1.count_dt\[4\] VGND VPWR
+ sky130_fd_sc_hd__or2b_1
X_0979_ VGND VPWR _0433_ _0436_ Shift_Register_Inst.data_out\[11\] net20 _0430_ _0435_
+ VGND VPWR sky130_fd_sc_hd__a2111o_1
X_0833_ VPWR VGND _0329_ Signal_Generator_2_0phase_inst.count\[1\] Signal_Generator_2_0phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__and2_1
X_0902_ Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_180phase_inst.count\[1\]
+ Signal_Generator_2_180phase_inst.count\[2\] _0380_ Signal_Generator_2_180phase_inst.count\[3\]
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31ai_1
XFILLER_0_43_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0764_ _0277_ Signal_Generator_1_90phase_inst.count\[0\] Signal_Generator_1_90phase_inst.count\[1\]
+ Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[3\]
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
X_0695_ VGND VPWR _0186_ _0225_ _0187_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_1316_ VPWR VGND Signal_Generator_1_90phase_inst.count\[3\] _0089_ _0024_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1178_ VGND VPWR _0541_ _0554_ _0555_ _0535_ VGND VPWR sky130_fd_sc_hd__o21ai_1
X_1247_ VPWR VGND _0612_ Dead_Time_Generator_inst_1.dt\[3\] _0609_ VGND VPWR sky130_fd_sc_hd__and2_1
X_1032_ VPWR VGND Signal_Generator_2_90phase_inst.count\[4\] _0463_ _0466_ _0464_
+ Signal_Generator_2_180phase_inst.count\[4\] _0465_ VGND VPWR sky130_fd_sc_hd__a221o_1
X_1101_ VPWR VGND _0516_ _0446_ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_33_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0747_ VPWR VGND _0264_ Signal_Generator_1_90phase_inst.count\[1\] VGND VPWR sky130_fd_sc_hd__inv_2
X_0816_ VGND VPWR _0316_ _0310_ _0315_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_16_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0678_ VGND VPWR _0146_ _0213_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_208 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_3__f_Dead_Time_Generator_inst_1.clk VGND VPWR clknet_0_Dead_Time_Generator_inst_1.clk
+ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1015_ VPWR VGND _0076_ _0450_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_30_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_185 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1280_ VGND VPWR net30 _0632_ _0513_ _0180_ VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_0_25_43 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0995_ VPWR VGND _0058_ _0448_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0780_ VPWR VGND _0007_ net44 VGND VPWR sky130_fd_sc_hd__inv_2
X_1332_ VPWR VGND Signal_Generator_1_270phase_inst.count\[5\] _0105_ _0019_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1263_ VGND VPWR _0581_ _0593_ _0175_ VGND VPWR sky130_fd_sc_hd__nor2_1
Xinput5 VGND VPWR net5 d1[2] VGND VPWR sky130_fd_sc_hd__buf_1
X_1194_ _0571_ Dead_Time_Generator_inst_1.count_dt\[4\] net27 VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0978_ VGND VPWR _0435_ _0431_ net15 _0434_ Shift_Register_Inst.data_out\[10\] VGND
+ VPWR sky130_fd_sc_hd__o211a_1
X_0832_ _0328_ Signal_Generator_2_0phase_inst.count\[5\] Signal_Generator_2_0phase_inst.count\[4\]
+ _0326_ _0327_ VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
X_0901_ VPWR VGND _0379_ _0370_ _0377_ _0037_ net51 VGND VPWR sky130_fd_sc_hd__a22o_1
X_0763_ VPWR VGND _0276_ _0266_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_11_125 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_147 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1315_ VPWR VGND Signal_Generator_1_90phase_inst.count\[2\] _0088_ _0023_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_0694_ VGND VPWR _0141_ _0224_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1177_ _0551_ _0552_ _0554_ _0553_ VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
X_1246_ VGND VPWR _0606_ _0608_ _0610_ _0611_ VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_0_33_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1031_ VGND VPWR _0465_ _0216_ _0214_ Signal_Generator_2_270phase_inst.count\[4\]
+ VGND VPWR sky130_fd_sc_hd__and3_1
X_1100_ VPWR VGND _0095_ _0515_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0746_ VGND VPWR _0263_ Signal_Generator_1_90phase_inst.count\[5\] Signal_Generator_1_90phase_inst.count\[4\]
+ _0261_ _0262_ VGND VPWR sky130_fd_sc_hd__o31a_2
X_0815_ VPWR VGND Signal_Generator_1_270phase_inst.count\[2\] _0315_ _0308_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0677_ VGND VPWR _0213_ _0211_ _0212_ _0182_ VGND VPWR sky130_fd_sc_hd__mux2_1
X_1229_ _0597_ _0598_ _0599_ _0561_ VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_30_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_103 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_147 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1014_ VPWR VGND _0450_ _0446_ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_12_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0729_ VPWR VGND Signal_Generator_1_0phase_inst.count\[2\] _0250_ _0243_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0994_ VPWR VGND _0057_ _0448_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_11_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1331_ VGND VPWR clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0018_ _0104_ Signal_Generator_1_270phase_inst.count\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
Xinput6 VGND VPWR net6 d1[3] VGND VPWR sky130_fd_sc_hd__buf_1
X_1193_ VPWR VGND _0570_ net39 _0567_ VGND VPWR sky130_fd_sc_hd__and2_1
X_1262_ VGND VPWR _0513_ net33 _0621_ _0174_ VGND VPWR sky130_fd_sc_hd__o21ba_1
XFILLER_0_46_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0977_ VGND VPWR _0434_ Shift_Register_Inst.data_out\[9\] net22 VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_9_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_248 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0900_ VGND VPWR _0379_ _0373_ _0378_ VGND VPWR sky130_fd_sc_hd__or2_1
XPHY_90 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0831_ VPWR VGND _0327_ Signal_Generator_2_0phase_inst.direction VGND VPWR sky130_fd_sc_hd__inv_2
X_0762_ VGND VPWR _0261_ _0275_ _0274_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_0693_ VGND VPWR _0224_ net1 _0223_ Shift_Register_Inst.data_out\[11\] VGND VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_159 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1314_ VPWR VGND Signal_Generator_1_90phase_inst.count\[1\] _0087_ _0022_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
Xclkbuf_0_Dead_Time_Generator_inst_1.clk VGND VPWR Dead_Time_Generator_inst_1.clk
+ clknet_0_Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_1176_ VGND VPWR _0553_ _0549_ _0550_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1245_ VGND VPWR _0609_ Dead_Time_Generator_inst_1.dt\[2\] _0607_ Dead_Time_Generator_inst_1.dt\[3\]
+ _0610_ VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_0_42_240 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1030_ _0464_ _0214_ _0216_ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
X_0814_ VPWR VGND Signal_Generator_1_270phase_inst.count\[2\] _0314_ _0311_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0745_ VPWR VGND _0262_ Signal_Generator_1_90phase_inst.direction VGND VPWR sky130_fd_sc_hd__inv_2
X_0676_ VGND VPWR _0186_ Shift_Register_Inst.shift_state\[2\] _0200_ _0212_ VGND VPWR
+ sky130_fd_sc_hd__or3b_1
X_1228_ VGND VPWR _0598_ Dead_Time_Generator_inst_2.count_dt\[1\] _0594_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_1159_ VGND VPWR _0536_ _0211_ _0208_ Signal_Generator_1_270phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_30_265 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_137 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_159 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1013_ VPWR VGND _0075_ _0449_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0728_ VPWR VGND Signal_Generator_1_0phase_inst.count\[2\] _0249_ _0246_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0659_ VGND VPWR _0151_ _0199_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_207 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_184 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_187 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0993_ VPWR VGND _0056_ _0448_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_1_221 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_168 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1330_ VGND VPWR clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0017_ _0103_ Signal_Generator_1_270phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1261_ VGND VPWR _0622_ _0621_ _0513_ _0173_ VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_0_36_99 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xinput7 VGND VPWR net7 d1[4] VGND VPWR sky130_fd_sc_hd__buf_1
X_1192_ VGND VPWR _0564_ _0566_ _0568_ _0569_ VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_0_46_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0976_ VPWR VGND _0433_ _0432_ net17 VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_0_13_190 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0830_ VPWR VGND Signal_Generator_2_0phase_inst.count\[1\] Signal_Generator_2_0phase_inst.count\[2\]
+ Signal_Generator_2_0phase_inst.count\[3\] Signal_Generator_2_0phase_inst.count\[0\]
+ _0326_ VGND VPWR sky130_fd_sc_hd__or4_2
XPHY_80 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0761_ Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[1\]
+ Signal_Generator_1_90phase_inst.count\[0\] _0274_ Signal_Generator_1_90phase_inst.count\[3\]
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31ai_1
X_0692_ _0187_ _0188_ _0223_ _0186_ VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
X_1313_ VPWR VGND Signal_Generator_1_90phase_inst.count\[0\] _0086_ _0021_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1244_ VPWR VGND _0609_ Dead_Time_Generator_inst_3.count_dt\[3\] VGND VPWR sky130_fd_sc_hd__inv_2
X_1175_ VPWR VGND _0548_ _0547_ _0542_ _0552_ VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_0_6_121 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0959_ VPWR VGND _0421_ Dead_Time_Generator_inst_1.go VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_17_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput10 VGND VPWR net10 d2[1] VGND VPWR sky130_fd_sc_hd__buf_1
X_0813_ VPWR VGND _0312_ _0020_ _0313_ _0015_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0744_ VPWR VGND Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[0\]
+ Signal_Generator_1_90phase_inst.count\[1\] Signal_Generator_1_90phase_inst.count\[3\]
+ _0261_ VGND VPWR sky130_fd_sc_hd__or4_2
X_0675_ VPWR VGND _0211_ Shift_Register_Inst.data_out\[6\] VGND VPWR sky130_fd_sc_hd__buf_2
X_1158_ VGND VPWR _0228_ _0530_ _0534_ _0535_ VGND VPWR sky130_fd_sc_hd__o21a_1
X_1227_ VGND VPWR _0597_ Dead_Time_Generator_inst_2.count_dt\[0\] Dead_Time_Generator_inst_2.count_dt\[1\]
+ _0593_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1089_ VPWR VGND _0085_ _0450_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1012_ VPWR VGND _0074_ _0449_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_12_200 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0727_ VPWR VGND _0247_ _0006_ _0248_ _0001_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0658_ VGND VPWR _0199_ Dead_Time_Generator_inst_1.dt\[1\] _0198_ _0182_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_230 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_199 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0992_ VPWR VGND _0448_ _0447_ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_41_103 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput8 VGND VPWR net8 d1[5] VGND VPWR sky130_fd_sc_hd__buf_1
X_1260_ VPWR VGND _0618_ Dead_Time_Generator_inst_3.count_dt\[2\] net45 _0622_ VGND
+ VPWR sky130_fd_sc_hd__a21oi_1
X_1191_ VGND VPWR _0567_ Dead_Time_Generator_inst_1.dt\[2\] _0565_ Dead_Time_Generator_inst_1.dt\[3\]
+ _0568_ VGND VPWR sky130_fd_sc_hd__o22a_1
X_0975_ VGND VPWR _0431_ Shift_Register_Inst.data_out\[10\] _0432_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_45_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_4__f_Dead_Time_Generator_inst_1.clk VGND VPWR clknet_0_Dead_Time_Generator_inst_1.clk
+ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
XPHY_81 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0760_ VPWR VGND _0273_ _0263_ _0271_ _0023_ net54 VGND VPWR sky130_fd_sc_hd__a22o_1
XPHY_92 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_25 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0691_ VGND VPWR _0142_ _0222_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1312_ VPWR VGND Signal_Generator_1_90phase_inst.direction _0085_ _0027_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1174_ VGND VPWR _0551_ _0548_ _0547_ _0542_ _0549_ _0550_ VGND VPWR sky130_fd_sc_hd__a32o_1
X_1243_ VPWR VGND Dead_Time_Generator_inst_1.dt\[2\] _0604_ Dead_Time_Generator_inst_1.dt\[1\]
+ _0608_ _0607_ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_19_228 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0889_ VPWR VGND _0371_ Signal_Generator_2_180phase_inst.count\[1\] Signal_Generator_2_180phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_0_42_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0958_ VGND VPWR net18 _0420_ VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_10_161 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput11 VGND VPWR net11 d2[2] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0743_ _0005_ _0244_ Signal_Generator_1_0phase_inst.direction Signal_Generator_1_0phase_inst.count\[4\]
+ _0260_ VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
X_0812_ VPWR VGND _0312_ _0307_ Signal_Generator_1_270phase_inst.direction _0313_
+ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0674_ VGND VPWR _0147_ _0210_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1157_ VGND VPWR _0533_ _0520_ Signal_Generator_1_0phase_inst.count\[1\] _0532_ _0534_
+ VGND VPWR sky130_fd_sc_hd__o22a_1
X_1226_ VGND VPWR _0164_ _0596_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1088_ VPWR VGND _0084_ _0450_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_2_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_212 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1011_ VPWR VGND _0073_ _0449_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0726_ VPWR VGND _0247_ _0242_ net58 _0248_ VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0657_ VPWR VGND _0194_ _0183_ Shift_Register_Inst.shift_state\[4\] _0198_ VGND VPWR
+ sky130_fd_sc_hd__or3_1
X_1209_ VGND VPWR net36 _0579_ _0581_ _0162_ VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_0_30_47 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_34 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_78 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_242 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0709_ VGND VPWR _0183_ Shift_Register_Inst.shift_state\[4\] Shift_Register_Inst.shift_state\[0\]
+ _0235_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_41_79 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0991_ VPWR VGND _0447_ _0446_ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_1_201 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_148 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_137 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1190_ VPWR VGND _0567_ Dead_Time_Generator_inst_1.count_dt\[3\] VGND VPWR sky130_fd_sc_hd__inv_2
Xinput9 VGND VPWR net9 d2[0] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_148 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0974_ VPWR VGND _0431_ Shift_Register_Inst.data_out\[9\] VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_45_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_82 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0690_ VGND VPWR _0222_ Shift_Register_Inst.data_out\[10\] _0221_ net1 VGND VPWR
+ sky130_fd_sc_hd__mux2_1
X_1311_ VGND VPWR clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0005_ _0084_ Signal_Generator_1_0phase_inst.count\[5\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1173_ VGND VPWR Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[2\]
+ Shift_Register_Inst.data_out\[5\] Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[2\]
+ _0211_ _0550_ VGND VPWR sky130_fd_sc_hd__mux4_1
X_1242_ VPWR VGND _0607_ Dead_Time_Generator_inst_3.count_dt\[2\] VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_27_251 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0888_ _0370_ Signal_Generator_2_180phase_inst.count\[5\] Signal_Generator_2_180phase_inst.count\[4\]
+ _0368_ _0369_ VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_42_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0957_ _0420_ _0413_ _0419_ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_0_10_173 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_240 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput12 VGND VPWR net12 d2[3] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0742_ _0260_ Signal_Generator_1_0phase_inst.count\[4\] Signal_Generator_1_0phase_inst.direction
+ _0240_ Signal_Generator_1_0phase_inst.count\[5\] VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
X_0673_ VGND VPWR _0210_ _0208_ _0209_ _0182_ VGND VPWR sky130_fd_sc_hd__mux2_1
X_0811_ VGND VPWR _0312_ _0311_ _0308_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1156_ VPWR VGND _0264_ _0208_ _0211_ _0533_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_1087_ VPWR VGND _0083_ _0450_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_28_6 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1225_ _0594_ _0595_ _0596_ _0561_ VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_30_224 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1010_ VPWR VGND _0072_ _0449_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_8_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_213 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0725_ VGND VPWR _0247_ _0246_ _0243_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0656_ VGND VPWR _0195_ _0152_ net60 VGND VPWR sky130_fd_sc_hd__xnor2_1
X_1208_ VPWR VGND _0559_ _0529_ _0558_ _0581_ _0560_ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_26_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1139_ VPWR VGND _0131_ _0447_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_7_240 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_176 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_46 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_59 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0708_ VGND VPWR _0137_ _0234_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0639_ VGND VPWR _0163_ _0185_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_190 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0990_ VGND VPWR net2 _0446_ VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_213 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_80 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0973_ VGND VPWR Shift_Register_Inst.data_out\[9\] Shift_Register_Inst.data_out\[10\]
+ _0430_ VGND VPWR sky130_fd_sc_hd__nor2_1
XPHY_83 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1310_ VGND VPWR clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0004_ _0083_ Signal_Generator_1_0phase_inst.count\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1241_ VGND VPWR _0606_ _0604_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_1.dt\[0\]
+ _0605_ VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_0_2_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1172_ VGND VPWR _0228_ _0549_ net5 VGND VPWR sky130_fd_sc_hd__or2b_1
XFILLER_0_27_263 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0956_ VGND VPWR _0419_ net3 _0228_ Dead_Time_Generator_inst_2.go VGND VPWR sky130_fd_sc_hd__mux2_1
X_0887_ VPWR VGND _0369_ Signal_Generator_2_180phase_inst.direction VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_33_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput13 VGND VPWR net13 d2[4] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0810_ VGND VPWR Signal_Generator_1_270phase_inst.count\[1\] Signal_Generator_1_270phase_inst.count\[0\]
+ _0311_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0741_ VGND VPWR _0004_ _0258_ _0257_ Signal_Generator_1_0phase_inst.direction _0242_
+ _0259_ VGND VPWR sky130_fd_sc_hd__a32o_1
X_0672_ VGND VPWR _0186_ Shift_Register_Inst.shift_state\[2\] _0196_ _0209_ VGND VPWR
+ sky130_fd_sc_hd__or3b_1
X_1224_ VGND VPWR _0595_ Dead_Time_Generator_inst_2.count_dt\[0\] _0593_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_1155_ _0532_ Signal_Generator_1_270phase_inst.count\[1\] _0211_ _0208_ _0531_ VGND
+ VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
X_1086_ VPWR VGND _0082_ _0450_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0939_ VGND VPWR _0046_ _0407_ _0406_ Signal_Generator_2_270phase_inst.direction
+ _0391_ _0408_ VGND VPWR sky130_fd_sc_hd__a32o_1
XFILLER_0_23_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_236 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_203 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_69 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_269 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0724_ VGND VPWR Signal_Generator_1_0phase_inst.count\[1\] Signal_Generator_1_0phase_inst.count\[0\]
+ _0246_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0655_ VGND VPWR _0196_ _0153_ _0197_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_1207_ VGND VPWR net41 _0579_ _0561_ _0161_ VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_0_19_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1069_ VPWR VGND _0501_ _0497_ _0502_ _0503_ VGND VPWR sky130_fd_sc_hd__a21o_1
X_1138_ VPWR VGND _0130_ _0447_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_7_252 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold2 VGND VPWR Dead_Time_Generator_inst_1.dt\[4\] net27 VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_0707_ VGND VPWR _0234_ net1 _0233_ net64 VGND VPWR sky130_fd_sc_hd__mux2_1
X_0638_ VGND VPWR _0185_ Dead_Time_Generator_inst_1.dt\[0\] _0184_ _0182_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_103 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_60 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0972_ VPWR VGND _0429_ Shift_Register_Inst.data_out\[12\] VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_42_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_84 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_62 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_51 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1171_ VGND VPWR _0548_ Signal_Generator_1_0phase_inst.count\[3\] _0520_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_1240_ VPWR VGND _0605_ Dead_Time_Generator_inst_3.count_dt\[0\] VGND VPWR sky130_fd_sc_hd__inv_2
X_0886_ VPWR VGND Signal_Generator_2_180phase_inst.count\[1\] Signal_Generator_2_180phase_inst.count\[2\]
+ Signal_Generator_2_180phase_inst.count\[3\] Signal_Generator_2_180phase_inst.count\[0\]
+ _0368_ VGND VPWR sky130_fd_sc_hd__or4_2
X_0955_ VPWR VGND net23 _0418_ VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
X_1369_ Dead_Time_Generator_inst_2.count_dt\[2\] clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
+ _0166_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput14 VGND VPWR net14 d2[5] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0740_ VGND VPWR _0240_ _0259_ Signal_Generator_1_0phase_inst.count\[4\] VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
X_0671_ VPWR VGND _0208_ Shift_Register_Inst.data_out\[5\] VGND VPWR sky130_fd_sc_hd__buf_2
X_1154_ Shift_Register_Inst.data_out\[5\] Shift_Register_Inst.data_out\[6\] _0531_
+ Signal_Generator_1_180phase_inst.count\[1\] VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
X_1223_ VPWR VGND _0594_ _0593_ Dead_Time_Generator_inst_2.count_dt\[0\] VGND VPWR
+ sky130_fd_sc_hd__and2_1
X_1085_ VPWR VGND _0081_ _0450_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0869_ VPWR VGND _0354_ _0055_ _0355_ _0050_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0938_ VGND VPWR _0389_ _0408_ Signal_Generator_2_270phase_inst.count\[4\] VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_215 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0723_ VPWR VGND _0000_ net42 VGND VPWR sky130_fd_sc_hd__inv_2
X_0654_ VGND VPWR _0194_ net57 _0197_ net48 VGND VPWR sky130_fd_sc_hd__o21ai_1
X_1206_ VPWR VGND _0576_ Dead_Time_Generator_inst_1.count_dt\[2\] net40 _0580_ VGND
+ VPWR sky130_fd_sc_hd__a21oi_1
X_1137_ VPWR VGND _0129_ _0447_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_7_264 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1068_ VPWR VGND _0502_ net10 VGND VPWR sky130_fd_sc_hd__inv_2
Xhold3 net28 _0614_ VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_0706_ VGND VPWR _0233_ _0187_ _0186_ _0188_ VGND VPWR sky130_fd_sc_hd__and3_1
Xclkbuf_3_5__f_Dead_Time_Generator_inst_1.clk VGND VPWR clknet_0_Dead_Time_Generator_inst_1.clk
+ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0637_ VPWR VGND Shift_Register_Inst.shift_state\[0\] _0183_ Shift_Register_Inst.shift_state\[4\]
+ _0184_ VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_0_35_159 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_83 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_50 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_129 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_192 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_140 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0971_ VGND VPWR net20 _0428_ VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_13_140 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_30 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_63 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1170_ VPWR VGND _0544_ _0546_ _0545_ _0543_ _0547_ VGND VPWR sky130_fd_sc_hd__or4_1
X_0885_ _0054_ _0351_ Signal_Generator_2_90phase_inst.direction Signal_Generator_2_90phase_inst.count\[4\]
+ _0367_ VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
X_0954_ VPWR VGND _0416_ _0417_ _0413_ _0418_ VGND VPWR sky130_fd_sc_hd__or3_1
X_1368_ Dead_Time_Generator_inst_2.count_dt\[1\] clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
+ _0165_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_1299_ VGND VPWR clknet_1_0__leaf_CLK_SR _0152_ _0073_ Shift_Register_Inst.shift_state\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0670_ VGND VPWR _0148_ _0207_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1084_ VPWR VGND _0080_ _0450_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1153_ VPWR VGND _0530_ net4 VGND VPWR sky130_fd_sc_hd__inv_2
X_1222_ _0593_ _0589_ _0590_ _0591_ _0592_ VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
X_0868_ VPWR VGND _0354_ _0349_ net52 _0355_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0799_ VGND VPWR _0285_ _0301_ _0302_ _0011_ _0303_ VGND VPWR sky130_fd_sc_hd__a2bb2o_1
X_0937_ VGND VPWR _0407_ Signal_Generator_2_270phase_inst.count\[4\] _0393_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_0722_ VGND VPWR _0242_ _0245_ _0006_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0653_ VGND VPWR _0194_ _0195_ Shift_Register_Inst.shift_state\[1\] _0196_ VGND VPWR
+ sky130_fd_sc_hd__or3_2
X_1067_ VPWR VGND _0498_ _0500_ _0499_ _0471_ _0501_ VGND VPWR sky130_fd_sc_hd__or4_1
X_1205_ VGND VPWR _0579_ Dead_Time_Generator_inst_1.count_dt\[2\] Dead_Time_Generator_inst_1.count_dt\[3\]
+ _0576_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1136_ VPWR VGND _0128_ _0447_ VGND VPWR sky130_fd_sc_hd__inv_2
Xhold4 net29 _0615_ VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0636_ VGND VPWR Shift_Register_Inst.shift_state\[2\] Shift_Register_Inst.shift_state\[1\]
+ Shift_Register_Inst.shift_state\[3\] _0183_ VGND VPWR sky130_fd_sc_hd__or3_2
X_0705_ VGND VPWR _0138_ _0232_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_94 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1119_ VPWR VGND _0112_ _0517_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_1_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_17 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_193 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0970_ VGND VPWR _0422_ _0428_ _0424_ VGND VPWR sky130_fd_sc_hd__or2b_1
X_1384_ Dead_Time_Generator_inst_3.go clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
+ _0181_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_60 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_233 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0884_ _0367_ Signal_Generator_2_90phase_inst.count\[4\] Signal_Generator_2_90phase_inst.direction
+ _0347_ Signal_Generator_2_90phase_inst.count\[5\] VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_12_74 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0953_ VGND VPWR _0228_ Dead_Time_Generator_inst_3.go _0417_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1367_ Dead_Time_Generator_inst_2.count_dt\[0\] clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
+ _0164_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_1298_ VGND VPWR clknet_1_0__leaf_CLK_SR _0151_ _0072_ Dead_Time_Generator_inst_1.dt\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_CLK_SR VGND VPWR clknet_0_CLK_SR clknet_1_1__leaf_CLK_SR VGND VPWR
+ sky130_fd_sc_hd__clkbuf_16
X_1221_ VGND VPWR net27 _0592_ Dead_Time_Generator_inst_2.count_dt\[4\] VGND VPWR
+ sky130_fd_sc_hd__or2b_1
X_1083_ VPWR VGND _0079_ _0450_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1152_ VGND VPWR _0525_ _0529_ _0528_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_0936_ VGND VPWR Signal_Generator_2_270phase_inst.count\[5\] Signal_Generator_2_270phase_inst.count\[4\]
+ _0403_ _0406_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_15_203 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0867_ VGND VPWR _0354_ _0353_ _0350_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0798_ VGND VPWR _0283_ _0303_ Signal_Generator_1_180phase_inst.count\[4\] VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_269 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0721_ VGND VPWR _0245_ Signal_Generator_1_0phase_inst.count\[4\] Signal_Generator_1_0phase_inst.count\[5\]
+ _0244_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0652_ VPWR VGND _0195_ _0183_ Shift_Register_Inst.shift_state\[4\] VGND VPWR sky130_fd_sc_hd__and2_1
X_1204_ VGND VPWR _0561_ _0578_ _0160_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_20_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_40 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1066_ VGND VPWR _0500_ _0216_ _0214_ Signal_Generator_2_270phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__and3_1
X_1135_ VPWR VGND _0127_ _0447_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0919_ VGND VPWR _0394_ Signal_Generator_2_270phase_inst.count\[4\] Signal_Generator_2_270phase_inst.count\[5\]
+ _0393_ VGND VPWR sky130_fd_sc_hd__and3_1
Xhold5 net30 Dead_Time_Generator_inst_4.count_dt\[4\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_125 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0635_ VPWR VGND _0182_ net1 VGND VPWR sky130_fd_sc_hd__buf_2
X_0704_ VGND VPWR _0232_ Shift_Register_Inst.data_out\[14\] _0231_ net1 VGND VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_71 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1049_ VGND VPWR _0483_ Signal_Generator_2_0phase_inst.count\[3\] _0467_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_1118_ VPWR VGND _0111_ _0517_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_34_150 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_131 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1383_ Dead_Time_Generator_inst_4.count_dt\[4\] clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
+ _0180_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_72 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_204 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0952_ VPWR VGND _0416_ net4 _0228_ VGND VPWR sky130_fd_sc_hd__and2_1
X_0883_ VGND VPWR _0053_ _0365_ _0364_ net52 _0349_ _0366_ VGND VPWR sky130_fd_sc_hd__a32o_1
XFILLER_0_12_97 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1366_ VGND VPWR clknet_1_0__leaf_CLK_SR _0163_ _0134_ Dead_Time_Generator_inst_1.dt\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1297_ VGND VPWR clknet_1_0__leaf_CLK_SR _0150_ _0071_ Dead_Time_Generator_inst_1.dt\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_270 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1151_ VPWR VGND _0526_ _0519_ _0524_ _0528_ _0527_ VGND VPWR sky130_fd_sc_hd__a22o_1
X_1220_ _0591_ Dead_Time_Generator_inst_2.count_dt\[4\] net27 VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__and2b_1
X_1082_ VPWR VGND _0078_ _0450_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0866_ VGND VPWR Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[1\]
+ _0353_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0935_ VPWR VGND _0405_ _0391_ _0402_ _0045_ Signal_Generator_2_270phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_15_215 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0797_ VGND VPWR _0287_ Signal_Generator_1_180phase_inst.direction _0302_ Signal_Generator_1_180phase_inst.count\[4\]
+ VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_62 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1349_ VPWR VGND Signal_Generator_2_180phase_inst.count\[1\] _0122_ _0036_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_0720_ VGND VPWR _0244_ Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[3\]
+ _0243_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0651_ VPWR VGND _0194_ Shift_Register_Inst.shift_state\[0\] VGND VPWR sky130_fd_sc_hd__inv_2
X_1134_ VPWR VGND _0126_ _0447_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1203_ VGND VPWR _0576_ _0578_ net63 VGND VPWR sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_52 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1065_ _0214_ _0216_ _0499_ Signal_Generator_2_180phase_inst.count\[1\] VGND VPWR
+ VGND VPWR sky130_fd_sc_hd__and3b_1
X_0849_ _0341_ Signal_Generator_2_0phase_inst.count\[2\] Signal_Generator_2_0phase_inst.count\[1\]
+ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[3\]
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
X_0918_ VGND VPWR _0393_ Signal_Generator_2_270phase_inst.count\[2\] Signal_Generator_2_270phase_inst.count\[3\]
+ _0392_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_11_251 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_137 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xhold6 net31 Dead_Time_Generator_inst_2.count_dt\[4\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_0703_ VGND VPWR _0231_ _0225_ _0200_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1117_ VPWR VGND _0110_ _0517_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_45_83 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_63 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1048_ VPWR VGND _0479_ _0481_ _0480_ _0471_ _0482_ VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_0_28_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_30 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_165 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_121 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1382_ Dead_Time_Generator_inst_4.count_dt\[3\] clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
+ _0179_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_11 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0882_ VGND VPWR _0347_ _0366_ Signal_Generator_2_90phase_inst.count\[4\] VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_216 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0951_ VGND VPWR net16 _0415_ VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_10_102 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1365_ Dead_Time_Generator_inst_1.count_dt\[4\] clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
+ _0162_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_1296_ VGND VPWR clknet_1_0__leaf_CLK_SR _0149_ _0070_ Dead_Time_Generator_inst_1.dt\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1150_ VGND VPWR Signal_Generator_1_90phase_inst.count\[4\] Signal_Generator_1_0phase_inst.count\[4\]
+ _0208_ Signal_Generator_1_270phase_inst.count\[4\] Signal_Generator_1_180phase_inst.count\[4\]
+ _0211_ _0527_ VGND VPWR sky130_fd_sc_hd__mux4_1
X_1081_ VGND VPWR _0157_ _0514_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0865_ VPWR VGND _0049_ net46 VGND VPWR sky130_fd_sc_hd__inv_2
X_0934_ VPWR VGND _0404_ _0403_ _0394_ _0405_ VGND VPWR sky130_fd_sc_hd__a21o_1
Xclkbuf_3_6__f_Dead_Time_Generator_inst_1.clk VGND VPWR net26 clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_238 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0796_ VGND VPWR _0301_ Signal_Generator_1_180phase_inst.count\[4\] _0300_ _0287_
+ VGND VPWR sky130_fd_sc_hd__and3_1
X_1348_ VPWR VGND Signal_Generator_2_180phase_inst.count\[0\] _0121_ _0035_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1279_ VGND VPWR _0179_ _0634_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0650_ VGND VPWR _0154_ _0193_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_241 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1064_ _0216_ Signal_Generator_2_90phase_inst.count\[1\] _0498_ _0214_ VGND VPWR
+ VGND VPWR sky130_fd_sc_hd__and3b_1
X_1133_ VPWR VGND _0125_ _0518_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1202_ VGND VPWR _0577_ _0576_ _0561_ _0159_ VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_0_18_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_64 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0848_ VPWR VGND _0340_ _0330_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0917_ VPWR VGND _0392_ Signal_Generator_2_270phase_inst.count\[1\] Signal_Generator_2_270phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__and2_1
X_0779_ VGND VPWR _0285_ _0288_ _0013_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_11_263 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_CLK_SR VGND VPWR CLK_SR clknet_0_CLK_SR VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xhold7 net32 Signal_Generator_2_270phase_inst.count\[0\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_0702_ VGND VPWR _0139_ _0230_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1116_ VPWR VGND _0109_ _0517_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1047_ VGND VPWR _0481_ Shift_Register_Inst.data_out\[8\] Shift_Register_Inst.data_out\[7\]
+ Signal_Generator_2_270phase_inst.count\[3\] VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_45_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_75 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_177 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1381_ Dead_Time_Generator_inst_4.count_dt\[2\] clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
+ _0178_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_149 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_236 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_67 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0881_ VGND VPWR _0365_ Signal_Generator_2_90phase_inst.count\[4\] _0351_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
XFILLER_0_12_55 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_228 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0950_ _0415_ _0413_ _0414_ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
X_1364_ Dead_Time_Generator_inst_1.count_dt\[3\] clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
+ _0161_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_1295_ VGND VPWR clknet_1_0__leaf_CLK_SR _0148_ _0069_ Dead_Time_Generator_inst_1.dt\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1080_ _0514_ _0461_ _0513_ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
X_0864_ VGND VPWR _0349_ _0352_ _0055_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0933_ _0404_ Signal_Generator_2_270phase_inst.count\[2\] Signal_Generator_2_270phase_inst.count\[1\]
+ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[3\]
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
X_0795_ VPWR VGND _0300_ Signal_Generator_1_180phase_inst.count\[5\] VGND VPWR sky130_fd_sc_hd__inv_2
X_1347_ VPWR VGND Signal_Generator_2_180phase_inst.direction _0120_ _0041_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1278_ _0632_ _0633_ _0634_ _0512_ VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
X_1201_ VGND VPWR net49 _0574_ _0577_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_20_253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1063_ VGND VPWR _0497_ Signal_Generator_2_0phase_inst.count\[1\] _0467_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_1132_ VPWR VGND _0124_ _0518_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0916_ _0391_ Signal_Generator_2_270phase_inst.count\[5\] Signal_Generator_2_270phase_inst.count\[4\]
+ _0389_ _0390_ VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
X_0847_ VGND VPWR _0326_ _0339_ _0338_ VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_0_11_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0778_ VGND VPWR _0288_ Signal_Generator_1_180phase_inst.count\[4\] Signal_Generator_1_180phase_inst.count\[5\]
+ _0287_ VGND VPWR sky130_fd_sc_hd__and3_1
Xhold8 net33 Dead_Time_Generator_inst_3.count_dt\[4\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_0701_ VGND VPWR _0230_ _0228_ _0229_ net1 VGND VPWR sky130_fd_sc_hd__mux2_1
X_1115_ VPWR VGND _0108_ _0517_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1046_ Shift_Register_Inst.data_out\[8\] Signal_Generator_2_90phase_inst.count\[3\]
+ _0480_ Shift_Register_Inst.data_out\[7\] VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_3_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_131 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_101 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1029_ _0463_ _0216_ _0214_ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
X_1380_ Dead_Time_Generator_inst_4.count_dt\[1\] clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
+ _0177_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_101 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_13 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_226 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_68 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_215 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0880_ VGND VPWR Signal_Generator_2_90phase_inst.count\[5\] Signal_Generator_2_90phase_inst.count\[4\]
+ _0361_ _0364_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_6_109 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1363_ Dead_Time_Generator_inst_1.count_dt\[2\] clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
+ _0160_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_1294_ VGND VPWR clknet_1_1__leaf_CLK_SR _0147_ _0068_ Shift_Register_Inst.data_out\[5\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_207 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0932_ VPWR VGND _0403_ _0393_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0863_ VGND VPWR _0352_ Signal_Generator_2_90phase_inst.count\[4\] Signal_Generator_2_90phase_inst.count\[5\]
+ _0351_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0794_ VPWR VGND _0299_ _0285_ _0296_ _0010_ net55 VGND VPWR sky130_fd_sc_hd__a22o_1
X_1346_ VGND VPWR clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0054_ _0119_ Signal_Generator_2_90phase_inst.count\[5\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1277_ _0633_ _0623_ Dead_Time_Generator_inst_4.count_dt\[1\] Dead_Time_Generator_inst_4.count_dt\[2\]
+ Dead_Time_Generator_inst_4.count_dt\[3\] VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_14_240 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1200_ VGND VPWR _0576_ Dead_Time_Generator_inst_1.count_dt\[0\] Dead_Time_Generator_inst_1.count_dt\[1\]
+ _0573_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1131_ VPWR VGND _0123_ _0518_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1062_ VGND VPWR Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[0\]
+ _0214_ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_180phase_inst.count\[0\]
+ _0216_ _0496_ VGND VPWR sky130_fd_sc_hd__mux4_1
XFILLER_0_34_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0915_ VPWR VGND _0390_ Signal_Generator_2_270phase_inst.direction VGND VPWR sky130_fd_sc_hd__inv_2
X_0846_ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[1\]
+ Signal_Generator_2_0phase_inst.count\[2\] _0338_ Signal_Generator_2_0phase_inst.count\[3\]
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31ai_1
X_0777_ VGND VPWR _0287_ Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[3\]
+ _0286_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_45_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1329_ VGND VPWR clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0016_ _0102_ Signal_Generator_1_270phase_inst.count\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_184 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold9 net34 Signal_Generator_2_0phase_inst.count\[0\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_218 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0700_ VGND VPWR _0229_ _0225_ _0196_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1114_ VPWR VGND _0107_ _0517_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_45_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_98 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1045_ Shift_Register_Inst.data_out\[7\] Shift_Register_Inst.data_out\[8\] _0479_
+ Signal_Generator_2_180phase_inst.count\[3\] VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_9_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0829_ _0019_ _0309_ Signal_Generator_1_270phase_inst.direction Signal_Generator_1_270phase_inst.count\[4\]
+ _0325_ VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_40_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_11 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_221 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_232 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1028_ VPWR VGND _0462_ net13 VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_16_165 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_14 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_216 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1293_ VGND VPWR clknet_1_1__leaf_CLK_SR _0146_ _0067_ Shift_Register_Inst.data_out\[6\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1362_ Dead_Time_Generator_inst_1.count_dt\[1\] clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk
+ _0159_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_227 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_230 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_271 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0862_ VGND VPWR _0351_ Signal_Generator_2_90phase_inst.count\[2\] Signal_Generator_2_90phase_inst.count\[3\]
+ _0350_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0931_ VGND VPWR _0389_ _0402_ _0401_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_0793_ VPWR VGND _0298_ _0297_ _0288_ _0299_ VGND VPWR sky130_fd_sc_hd__a21o_1
Xrebuffer1 VGND VPWR clknet_0_Dead_Time_Generator_inst_1.clk net26 VGND VPWR sky130_fd_sc_hd__buf_8
X_1345_ VPWR VGND Signal_Generator_2_90phase_inst.count\[4\] _0118_ _0053_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_1276_ VGND VPWR _0632_ Dead_Time_Generator_inst_4.count_dt\[2\] Dead_Time_Generator_inst_4.count_dt\[3\]
+ _0626_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1130_ VPWR VGND _0122_ _0518_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_7_205 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1061_ VPWR VGND _0495_ net9 VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_34_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0845_ VPWR VGND _0337_ _0328_ _0335_ _0030_ net69 VGND VPWR sky130_fd_sc_hd__a22o_1
X_0914_ VPWR VGND Signal_Generator_2_270phase_inst.count\[1\] Signal_Generator_2_270phase_inst.count\[2\]
+ Signal_Generator_2_270phase_inst.count\[3\] Signal_Generator_2_270phase_inst.count\[0\]
+ _0389_ VGND VPWR sky130_fd_sc_hd__or4_2
X_0776_ VPWR VGND _0286_ Signal_Generator_1_180phase_inst.count\[0\] Signal_Generator_1_180phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_0_38_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1328_ VGND VPWR clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0015_ _0101_ Signal_Generator_1_270phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1259_ VGND VPWR _0621_ Dead_Time_Generator_inst_3.count_dt\[2\] Dead_Time_Generator_inst_3.count_dt\[3\]
+ _0618_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_46_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1113_ VPWR VGND _0106_ _0517_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1044_ VPWR VGND _0478_ net12 VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_10_90 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0759_ VGND VPWR _0273_ _0267_ _0272_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0828_ _0325_ Signal_Generator_1_270phase_inst.count\[4\] Signal_Generator_1_270phase_inst.direction
+ _0305_ Signal_Generator_1_270phase_inst.count\[5\] VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_40_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_244 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1027_ _0461_ _0457_ _0458_ _0459_ _0460_ VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_16_177 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_7__f_Dead_Time_Generator_inst_1.clk VGND VPWR net26 clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_44 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_206 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_191 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_14 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_36 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_239 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1361_ Dead_Time_Generator_inst_1.count_dt\[0\] clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk
+ _0158_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_1292_ VGND VPWR clknet_1_0__leaf_CLK_SR _0145_ _0066_ Shift_Register_Inst.data_out\[7\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_155 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_242 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_46 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0861_ VPWR VGND _0350_ Signal_Generator_2_90phase_inst.count\[1\] Signal_Generator_2_90phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__and2_1
X_0930_ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[1\]
+ Signal_Generator_2_270phase_inst.count\[2\] _0401_ Signal_Generator_2_270phase_inst.count\[3\]
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31ai_1
X_0792_ _0298_ Signal_Generator_1_180phase_inst.count\[0\] Signal_Generator_1_180phase_inst.count\[1\]
+ Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[3\]
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_23_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1344_ VPWR VGND Signal_Generator_2_90phase_inst.count\[3\] _0117_ _0052_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1275_ VGND VPWR _0178_ _0631_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1060_ VPWR VGND _0491_ _0493_ _0492_ _0484_ _0494_ VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_0_7_228 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0844_ VGND VPWR _0337_ _0331_ _0336_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0913_ _0040_ _0372_ net68 Signal_Generator_2_180phase_inst.count\[4\] _0388_ VGND
+ VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
X_0775_ VGND VPWR _0285_ Signal_Generator_1_180phase_inst.count\[5\] Signal_Generator_1_180phase_inst.count\[4\]
+ _0283_ _0284_ VGND VPWR sky130_fd_sc_hd__o31a_2
X_1327_ VGND VPWR clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0014_ _0100_ Signal_Generator_1_270phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1258_ VGND VPWR _0513_ _0620_ _0172_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1189_ VPWR VGND Dead_Time_Generator_inst_1.dt\[2\] _0562_ Dead_Time_Generator_inst_1.dt\[1\]
+ _0566_ _0565_ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_46_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_34 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1043_ VGND VPWR _0475_ _0476_ _0469_ _0477_ VGND VPWR sky130_fd_sc_hd__or3b_1
X_1112_ VPWR VGND _0517_ _0446_ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_28_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_186 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0758_ VPWR VGND Signal_Generator_1_90phase_inst.count\[2\] _0272_ _0265_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0827_ VGND VPWR _0018_ _0323_ _0322_ Signal_Generator_1_270phase_inst.direction
+ _0307_ _0324_ VGND VPWR sky130_fd_sc_hd__a32o_1
X_0689_ VGND VPWR _0200_ Shift_Register_Inst.shift_state\[3\] Shift_Register_Inst.shift_state\[2\]
+ _0221_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_19_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_137 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1026_ VGND VPWR Dead_Time_Generator_inst_1.dt\[4\] _0460_ Dead_Time_Generator_inst_4.count_dt\[4\]
+ VGND VPWR sky130_fd_sc_hd__or2b_1
XFILLER_0_39_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_16 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1009_ VPWR VGND _0071_ _0449_ VGND VPWR sky130_fd_sc_hd__inv_2
XPHY_27 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_6 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1360_ VPWR VGND Signal_Generator_2_270phase_inst.count\[5\] _0133_ _0047_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1291_ VGND VPWR clknet_1_0__leaf_CLK_SR _0144_ _0065_ Shift_Register_Inst.data_out\[8\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0860_ VGND VPWR _0349_ Signal_Generator_2_90phase_inst.count\[5\] Signal_Generator_2_90phase_inst.count\[4\]
+ _0347_ _0348_ VGND VPWR sky130_fd_sc_hd__o31a_2
X_0791_ VPWR VGND _0297_ _0287_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1343_ VPWR VGND Signal_Generator_2_90phase_inst.count\[2\] _0116_ _0051_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_1274_ VGND VPWR _0631_ _0629_ _0513_ _0630_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0989_ VGND VPWR net25 _0445_ _0436_ _0429_ _0440_ VGND VPWR sky130_fd_sc_hd__a31o_4
X_0912_ _0388_ Signal_Generator_2_180phase_inst.count\[4\] Signal_Generator_2_180phase_inst.direction
+ _0368_ Signal_Generator_2_180phase_inst.count\[5\] VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
X_0843_ VPWR VGND Signal_Generator_2_0phase_inst.count\[2\] _0336_ _0329_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0774_ VPWR VGND _0284_ Signal_Generator_1_180phase_inst.direction VGND VPWR sky130_fd_sc_hd__inv_2
X_1326_ VGND VPWR clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0020_ _0099_ Signal_Generator_1_270phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1257_ VGND VPWR _0618_ _0620_ net62 VGND VPWR sky130_fd_sc_hd__xnor2_1
X_1188_ VPWR VGND _0565_ Dead_Time_Generator_inst_1.count_dt\[2\] VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_46_165 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_46 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1042_ VGND VPWR _0476_ _0470_ _0474_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_45_45 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1111_ VPWR VGND _0105_ _0516_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_43_102 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0757_ VPWR VGND Signal_Generator_1_90phase_inst.count\[2\] _0271_ _0268_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0826_ VGND VPWR _0305_ _0324_ Signal_Generator_1_270phase_inst.count\[4\] VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
X_0688_ VGND VPWR _0143_ _0220_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1309_ VGND VPWR clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0003_ _0082_ Signal_Generator_1_0phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_102 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_198 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1025_ _0459_ Dead_Time_Generator_inst_4.count_dt\[4\] Dead_Time_Generator_inst_1.dt\[4\]
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
X_0809_ VPWR VGND _0014_ net35 VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_31_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_205 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_68 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_116 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_17 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1008_ VPWR VGND _0070_ _0449_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_12_160 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1290_ VGND VPWR clknet_1_1__leaf_CLK_SR _0143_ _0064_ Shift_Register_Inst.data_out\[9\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_263 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_26 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0790_ VGND VPWR _0283_ _0296_ _0295_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_1342_ VPWR VGND Signal_Generator_2_90phase_inst.count\[1\] _0115_ _0050_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1273_ VGND VPWR _0630_ Dead_Time_Generator_inst_4.count_dt\[2\] _0626_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_0988_ VGND VPWR _0445_ _0444_ Shift_Register_Inst.data_out\[10\] _0431_ _0442_ VGND
+ VPWR sky130_fd_sc_hd__a31o_4
X_0842_ VPWR VGND Signal_Generator_2_0phase_inst.count\[2\] _0335_ _0332_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0911_ VGND VPWR _0039_ _0386_ _0385_ net51 _0370_ _0387_ VGND VPWR sky130_fd_sc_hd__a32o_1
XFILLER_0_11_225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0773_ VPWR VGND Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[0\]
+ Signal_Generator_1_180phase_inst.count\[1\] Signal_Generator_1_180phase_inst.count\[3\]
+ _0283_ VGND VPWR sky130_fd_sc_hd__or4_2
X_1325_ VPWR VGND Signal_Generator_1_180phase_inst.count\[5\] _0098_ _0012_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1256_ VGND VPWR _0619_ _0618_ _0513_ _0171_ VGND VPWR sky130_fd_sc_hd__nor3_1
X_1187_ VGND VPWR _0564_ _0562_ Dead_Time_Generator_inst_1.dt\[1\] _0563_ Dead_Time_Generator_inst_1.dt\[0\]
+ VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_0_6_241 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1110_ VPWR VGND _0104_ _0516_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_29_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1041_ VPWR VGND _0468_ _0470_ _0474_ _0475_ _0462_ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_9_57 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0825_ VGND VPWR _0323_ Signal_Generator_1_270phase_inst.count\[4\] _0309_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_0756_ VPWR VGND _0269_ _0027_ _0270_ _0022_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0687_ VGND VPWR _0220_ Shift_Register_Inst.data_out\[9\] _0219_ _0182_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
X_1308_ VGND VPWR clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0002_ _0081_ Signal_Generator_1_0phase_inst.count\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1239_ VPWR VGND _0604_ Dead_Time_Generator_inst_3.count_dt\[1\] VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_34_114 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_177 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1024_ _0458_ Dead_Time_Generator_inst_4.count_dt\[3\] Dead_Time_Generator_inst_1.dt\[3\]
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
X_0808_ VGND VPWR _0307_ _0310_ _0020_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0739_ VGND VPWR _0258_ Signal_Generator_1_0phase_inst.count\[4\] _0244_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
XFILLER_0_39_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_106 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_48 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_128 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_CLK_SR VGND VPWR clknet_0_CLK_SR clknet_1_0__leaf_CLK_SR VGND VPWR
+ sky130_fd_sc_hd__clkbuf_16
X_1007_ VPWR VGND _0069_ _0449_ VGND VPWR sky130_fd_sc_hd__inv_2
XPHY_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_220 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_212 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_38 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1341_ VPWR VGND Signal_Generator_2_90phase_inst.count\[0\] _0114_ _0049_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1272_ VGND VPWR Dead_Time_Generator_inst_4.count_dt\[2\] _0629_ _0626_ VGND VPWR
+ sky130_fd_sc_hd__nand2_1
X_0987_ VGND VPWR _0444_ Shift_Register_Inst.data_out\[12\] _0439_ _0443_ VGND VPWR
+ sky130_fd_sc_hd__and3_1
XFILLER_0_9_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0841_ VPWR VGND _0333_ _0034_ _0334_ _0029_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0910_ VGND VPWR _0368_ _0387_ Signal_Generator_2_180phase_inst.count\[4\] VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
X_0772_ _0026_ _0266_ Signal_Generator_1_90phase_inst.direction Signal_Generator_1_90phase_inst.count\[4\]
+ _0282_ VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
X_1324_ VPWR VGND Signal_Generator_1_180phase_inst.count\[4\] _0097_ _0011_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_1255_ VGND VPWR net50 _0616_ _0619_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1186_ VPWR VGND _0563_ Dead_Time_Generator_inst_1.count_dt\[0\] VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_6_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1040_ VGND VPWR _0473_ _0467_ Signal_Generator_2_0phase_inst.count\[5\] _0472_ _0474_
+ VGND VPWR sky130_fd_sc_hd__o22a_1
X_0755_ VPWR VGND _0269_ _0263_ net54 _0270_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0824_ VGND VPWR Signal_Generator_1_270phase_inst.count\[5\] Signal_Generator_1_270phase_inst.count\[4\]
+ _0319_ _0322_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_28_178 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0686_ VGND VPWR _0196_ Shift_Register_Inst.shift_state\[3\] _0187_ _0219_ VGND VPWR
+ sky130_fd_sc_hd__or3b_1
X_1169_ Shift_Register_Inst.data_out\[6\] Signal_Generator_1_90phase_inst.count\[3\]
+ _0546_ Shift_Register_Inst.data_out\[5\] VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_1
X_1307_ VGND VPWR clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0001_ _0080_ Signal_Generator_1_0phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_91 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1238_ VGND VPWR _0561_ _0573_ _0169_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1023_ VGND VPWR _0454_ _0455_ Dead_Time_Generator_inst_1.dt\[2\] _0451_ _0457_ _0456_
+ VGND VPWR sky130_fd_sc_hd__o221a_1
X_0738_ VGND VPWR Signal_Generator_1_0phase_inst.count\[5\] Signal_Generator_1_0phase_inst.count\[4\]
+ _0254_ _0257_ VGND VPWR sky130_fd_sc_hd__or3b_1
X_0807_ VGND VPWR _0310_ Signal_Generator_1_270phase_inst.count\[4\] Signal_Generator_1_270phase_inst.count\[5\]
+ _0309_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0669_ VGND VPWR _0207_ Dead_Time_Generator_inst_1.dt\[4\] _0206_ _0182_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_19 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1006_ VPWR VGND _0068_ _0449_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_16_93 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_232 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_126 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_246 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_118 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1340_ VPWR VGND Signal_Generator_2_90phase_inst.direction _0113_ _0055_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1271_ VGND VPWR _0177_ _0628_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0986_ VPWR VGND _0432_ net24 _0430_ _0443_ net19 VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_1_151 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0840_ VPWR VGND _0333_ _0328_ net59 _0334_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0771_ _0282_ Signal_Generator_1_90phase_inst.count\[4\] Signal_Generator_1_90phase_inst.direction
+ _0261_ Signal_Generator_1_90phase_inst.count\[5\] VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
X_1323_ VPWR VGND Signal_Generator_1_180phase_inst.count\[3\] _0096_ _0010_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1254_ VGND VPWR _0618_ Dead_Time_Generator_inst_3.count_dt\[0\] Dead_Time_Generator_inst_3.count_dt\[1\]
+ _0615_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1185_ VPWR VGND _0562_ Dead_Time_Generator_inst_1.count_dt\[1\] VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_46_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0969_ VGND VPWR net17 _0427_ VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_45_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0754_ VGND VPWR _0269_ _0268_ _0265_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0823_ VPWR VGND _0321_ _0307_ _0318_ _0017_ net61 VGND VPWR sky130_fd_sc_hd__a22o_1
X_0685_ VGND VPWR _0144_ _0218_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1306_ VGND VPWR clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0000_ _0079_ Signal_Generator_1_0phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1099_ VPWR VGND _0094_ _0515_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1168_ VGND VPWR _0545_ Shift_Register_Inst.data_out\[6\] Shift_Register_Inst.data_out\[5\]
+ Signal_Generator_1_270phase_inst.count\[3\] VGND VPWR sky130_fd_sc_hd__and3_1
X_1237_ VGND VPWR net31 _0601_ _0561_ _0168_ VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_0_42_171 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1022_ VGND VPWR Dead_Time_Generator_inst_1.dt\[3\] _0456_ Dead_Time_Generator_inst_4.count_dt\[3\]
+ VGND VPWR sky130_fd_sc_hd__or2b_1
X_0737_ VPWR VGND _0256_ _0242_ _0253_ _0003_ Signal_Generator_1_0phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__a22o_1
X_0806_ VGND VPWR _0309_ Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[3\]
+ _0308_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0668_ VGND VPWR _0186_ Shift_Register_Inst.shift_state\[2\] _0205_ _0206_ VGND VPWR
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_21_83 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_193 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xhold40 net65 Signal_Generator_2_0phase_inst.count\[4\] VGND VPWR VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_1005_ VPWR VGND _0067_ _0449_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_44_244 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_211 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_258 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_211 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
.ends

